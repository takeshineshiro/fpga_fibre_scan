��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	��q5.A��|�H����VM.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y_�L_H��-..i=?�m��+�<4��ˌ��|��v��ӳ��$Fe@���N�w	*D���y&�f��+K��[y��ڂ�Vs>�+��T�,F���J�/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&�z(ݲm@�)yH�I@'�ew2�\�蝆�u����l�|���j����1�}�<RK��2Ee�Y�R2
�I.��	���
�Ɛ��BR�[_i����v H�$�Yo�1z�:맷�m��d�78�^f��G�n�QX�v����<.���+��T���jB�Fg�:S�Q�[�$A�������6��H4�
� �AH�T�t��3��'�Wا[~�l]ǜ�����] ��F@�4%���D�Pfc����2P����/�"��< ���X�M+��tc��P9P��`�.�D���J7"� $��|�M
r:�����u��w)�S �J���vy7��Mv�9�E���5�n�Gb�Șo8�:r&@1�+Q�<Ǵoe� 2m�!=�y����h�}�)�����=nAIZ(�2��o?�M��;]\V�A}��}���V���8e3Z}�ax�� 5�k�8���҆�|n����vJ�^�R�!�"s�x��`x)J�Й�m�BdP*4�h־�-9�,����"��yА���kc�.[K��mN,����0j Oag�ì���Tl��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcz��9�L�*8h
����;�3.-D)>ƾ~���($�N��$�`���PЯ*{��i@F��X���I��`%�W8��6~ă��H>:벡^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�YZY0@ìOJ����%@����BF+�va��2鍔�	g\A^��+o��	g�yߓ����<�m��+��$|��;D���J7"�~�#�B7vC/��&)Y�{��n���Yk"1/�<4��ˌ��|��v���k.!�l�	�/�No`g	�ts�q�)3[�u8�����$G�yد�9�����~�����wl��h�)H��!n�'�\�J׽Z�ݽ;.p�7:SW�<�6�Q=Ի�弳$�.����~���kR$�kn���5���k�����L9��DUR�ߟ�;�Æ�MYi=�/M��%�p@Y�4Eb��ޒ`��`$���g>넽� �\Yy��M��(�K����!�ʭwV~���Vr�{r�����-N�'E�HG�vz��RxX��TԘ�H <8�k[p�M����G��u�c��Q��ݭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3j���T������q��
�e�~w�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�>.��̡��@��܊_�1���r�.v���t��W2�7�t`\���~��;�,!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�&�7m�3�i�V��wvf��q�d� s�\{]���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�z�-�v�k[�~�Z1~�g]�c�u��QF�s�����?!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD��� �oݗ����[2$L�e�(��0���N���z[�M�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD� ��*2�fNY��'�T��@�ш�ň6���D)9W �v:ι�Y7���&�_k�c��`�)\��FCR��]��e܅����
@{���e����q����؍��R��{QgkS�(!�`�(i3��%<�d�6�.�)��:�����y��j��k�s5=Ύ�9�j���B���7�F�ĭW�.�%6�<]"�:sNcbp��'�����U��ݚ�Н�`���*1R����
wL<65���Yl���#Kv���:1�#����az�~��c�&ck��K6�L+�.8%�����dN�<@Iv���a_|����ݚ�Н�H/�I��(B&�2�>��}YY�{'%s�&�
�0�pD��ZOU�g��U-�ee�@Rv����my$�N��o�/���;��6���m�XQ���z�+ N���>S̮�K�+EC�hHc�Ì49�����x�����s��l|�*"k���(ӈ��z&��)Q��!�`�(i3-Gb��F��E����Fv�Z��P,N�:2QYeƈ)P<�ܓ�Y���aR�!�`�(i3⤵�6�)�T<9 =��9�j���B�<Vo�eo���9�r7�K6�L+�.8%�����dN�<@Iv���a_|����ݚ�Н�ʅ|7@J=�P�:SôHaKv���ft�s� uƍ2���l�`���*1�I���`�����-VL�1���o�l����4�n���xǊj�ë��&�E���Kt�������qϛ�M~�ˇ�h��]�Hlu�����}Dq�f��H	EJF�dʀ�����
t��f"�	-7��8�r�%�
���lC��U7�C��zC@�D+���4Yq(����(p���	��
�Q�}A�����2�[<�!�� �w�;>cbp��'�����C��ݚ�Н��:#�R_��+�
�c�~��G1��[���J���T���b+}y[���S�fp�*x�$�Z�YBQ.K��]�!���\B��V���|e"h�wֈ�WI��}f����y���29��:|[%.�m�QA�Q* !�`�(i3H���L@�B�/�@TP3C6�HaDl����/	e�Ҏ�R]����pz�b'�tN2s���(����5��x���|�:S�Q�[����g��.�V�k�J8U��C�V�8��ݾ�]9!s�(����5��x���|�:S�Q�[����g��x�48<?���G-�43�J͇Z6W.d��N((�}���cbp��'��Q>��k���D�s�,7���a�W��l����4�n���xǊ�Ru�A^H�X~L��U��0���g�-�:���9�^���N�j�<�_�l����4�x�ߴ�2�rP���(�U�w�Q�q�v��:�����`�@��i���e�g5�<���e9�j���B���W�Ħ�〧I��ɳE��׆��d�٣���,�JL��ކ�|u�S
$�0�Q��v1a{J�_�S�
utY�{'%s���'����+D���0�7a
��r�"j���b7Z�n��[��{_8�Y��=�}�Vݨ���,D��9=Sr���n��a� _�S�
utY�{'%s�Ǹ2���;�¬pX��g��U-�ee�@Rv����my$�N�����X8��$��Xo���v&�7W�U�����}8���uӜk��(���B����ѾJJ�� ��˽��r�g��gQ�qs�r�hz7���&�_0M�/�s���Z�>)���'vX[��7�t`\�� ðc4u���0@ȹ��ZBi�mR�5*%ol��H�)g��i3�|)sՀ@���l�}�p��g��Bڎ@L�xg`�H�4��`t�A~�@����gG8���� 3��~᩷�������fG��G�62��`t�A~���	wD�B�щ%��� ���V�8�|���$���!<.S��!���d.W>	����h4!��a=�����`+iYbú��g�=�R��T�55��2@���G�>�o�5��ˇ���<�6�Q=�܇�7��:1|%�Ӿ�`^X�k��D���z����y��lDp��.^	O:�i�Eg�[`�f��$��|o����;���'T���+���\�]�2	�� �UI�����d��i��7�����h�ura$�>�Q�ˤK0���O잢+K�Bu~]�u;Q��5��Hf�v!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��FRv"(�����d�������r����!�`�(i3!�`�(i3!�`�(i3!�`�(i3�XW�����;��`�x�M�}�P��>������ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i36�e�:r�"2�?��4x.�bI	\������ˊ%<.�cs��'�)a��p�����x(�i��/R<��}�u�4���������]:��b�wi��Ȱ�(�φ��<�6������~�c!���d.W>	����hs�à���~���=�q1tSjv�!�`�(i3�LD��B����Y� ���Ja�~'T.,����/9�=e��n�_��&�(���D'?��uy���V���%g��Un��Pxκ�ǣ��ԩO�j���Gp��ܐ�}�г*O�v��b�*���]k�WM��q�U��)��N�2 �3�]�7�"�Ͻg�iO��|��h��èV8�w��U�Mg�w�u�$�&�V(*�O�qM�4�<>�[!�`�(i3�=0Zcs�ݚ�Н����v�gY�ڰ݉ �%��v��!�`�(i3�ݚ�Н��˸�կ���/8����_�mS8<�n�ݚ�Н�1���/���6�<"��
8�	3��Ra])n#���r����
��X��F��[�i�[e}��T�W���%>�rGO�D mWNG�&ց�*��W�"v�Q!�`�(i3o�;�6���|e"h�wֈ�WI��}f���#�+#��]ž_�F�i#\��u�F�;��ko_�mS8<�n�ݚ�Н�1���/������E�EczUEg�>
�:qEp'{w#/ B���S�f������f���5n��}Dq�f���Ě���ž_�Fȋ�O�������ϒ!�`�(i3��򴏓�	k	䶙%A��ʺ�l�?�{�XԔ�Z?�߸��S�Ȍ�l
�VD����-��Tc��փ6�o8:4��V���%��c�+5L{y����i�q,?5q�Y�ڒ���
�a(M���8���Q�t�vz�	�o���Ȋx��7��A0ɷ��9)P<�ܓ�Y-�E��%����I��毘3)�:i#\��u��.d�i�>1tSjv�c�@���Pxκ�ǣ���Y� �����"���jVѭ@P#+_]ݱ��3,l5�k	䶙%�F�}қ~���Ě�����[�"��$Q�s#�����>e-Gb��F�n��뾦�`
 ֢���V�ܔ�s
���NM���t�td���5l��5��\zm�$�ܻ�u��r��'E>����������f���5n��}Dq�f�1���~c�@���Pxκ�ǣ���Y� �>���������F��O�!�`�(i3N� ����V(pyL0D�!#��MP�3,l5�k	䶙%A��ʺ�l���4�CD5����+Y��a�U�ے
�,�j�<[�k]m���Ϩ�@k�,+��Z>³��$���!<.S�����*V�	m�]�� �k���L��?8��Cd[Uu��r��m����'K�j��=��\�{_8�Y��=�}�Vݨ�R� v+0x%�kˣ���3�|* ���dN�<@Iv��nt=:ྻ�!����.P�:�����3&�.C������٫Np�&�U��f���Aڬ&W�n�>oSbT��;�k��-�����
�*�ݡK�+���w�x~Pj.
��S�CП����S�f%�kˣ���3�|* ���Mp0բ����g��HN��R���ء�I�Ǡ�����߸��S�Ȍ��vZ��4-�k]m��4E������k]m���#�')�~=�yۂ�J1Cw�Hm���ǽbI��#��$���S~d6:��ft�� �yۂ�J1��S����D� �B��=��/ 0;��5,�O[p8�]�1����W� �EA��i.� �#�i���U]�%N\�*�q &��)f=L��#� �+=]�-S��\Ys|��yW��(�`n�>]˕�8�3�M)h�~������1;[lz!z1��,�gq� �ɰ5�*�"��y������6~0��R��4J���g?mЛR>l'�J<!��޳?%*3)t�O9�T�}���e��r�Ө/a�]v�����7}Wo�����:.e�^����pq5H(R�XY�kn�j��x߆�V�$
Ɏ�/��>3�%9���D��z�1�'싯��xQ17�b�����d���!iH/�I��(��"Jk�\K7͍��ճ��)��{��&^8��a�����y�w�a���Bƌ���� ���B�#9ʿT�;��|B <�Az��0�-GS'�i�*ڶ�UKs,���́m��BK�+���w�X�{̡�Z7���&�_��lC��U�T���rJ|�6soi���{r����r�gKG�͎F�c�|��J�C�CW�w��fDcW�b����w��-��Xo�H!.� �#�imWᅫw�5�O�%E#P�i����|M�U��b�z'hۉ)��ԩ�c!6j�"Hs��=��Ln�ŭ�s�=�Q��X�w��8�3�M�oT��O?�d���&��6)��Tj�`����nm����'KN+?��T�{r��;�¬pX��g��U-�e���O�s?�d���&��l��"q����Sv�Q{u�D�$�R����b