��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag������T-ǋ 4�i� ������[���a�8%`��4�s�6�XAoeuxLZ�#8v��fT��ı��¥���hM�,=i�@x_\q�jB�Fg�Y씤`��p��>�B�㬊�N�����3��>�U���T���딣0&_���X0���2|	p��rw@	@us��Nิi'Y0ii^sZ��yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��:K����HJ{D�9h�@dw.+��CS�����L�;���xI+r�� 0�D�A�f�mX��)D�b@��Ó���K^�7��5p�v�r�:�u)�~�<��[�T�٥��T���BR�[_ň��h��Ev�i<l��]a�{ڬ��;�Ӏ��nrm؊(�{�P�1|�+=ύ�-�����!Jė/�Ҏ/��?��\�D�PKA[[Nyx���GlVҤ�ן2#a����+�jԪ�"��)�k�5��i��$�Ƣ�/몍N�������=�����(��h�]X.�H@f�foS�EjLP� #V�r�O��C��0����"g�����I����oi21���fѶ^��7C��H�K��wAG6�i��<&����P'o#�D�Z�ǝ��RL�a)=�y�~ ���H7����En��"ydO�A�Eh�7C��H���j�v�?�]E�]�����+�ڔހ��g�R��b�^��\�}w�*
� �AH���g���	�e��ME
v���Fw4�Š�@`��F@�4%�?$7��fǜ��ǽ��"�-�vF�..���}�<�����_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢS����E@�gh1���Yh�\��q��r����N{a�9Ow�Y��k��ı��*���q{?d']l�f��Wj gs����'v�]wɭ�7��r�=!�`�(i3N�By3��<�]�!����M[��Ǣ)�k�4�U!�`�(i3�����5	���]����,�JL����?D�8��R�����!�`�(i3�����5	���]���>����CΌh��eZ!�`�(i3Y%T��BPe.��xu	�>��l%i�-�5`z��s�Ƀ�?PA�':E����j���0z�cUL�I��6���T�\ ��:E��]��8S�n�(�a�x�f7﹏N�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�����5	���]���>����CηxmQ,ۘS!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FH=Y��@�E����F7G#+��\w��0]�o�t��F�e{iʖ.	��A���TD��ό���.Ӂ��̰�!i�q8�2t�ݡ��1����(�
t��Y�{'%s2�ew�a(􆿳����^���(R\֎u�,��7-�)�V�3j@IE�U��>��l%i�-�jo�'q�!�`�(i3�E����F7G#+����w�V�"�"��FX1�������Pc��q�Pe:[e��m�D��L���_�L�Ȳ�V�溜��D�,�H�.�z,y������Ls�F�%ܪ���P}|��XH��/gt׶�h��y�xv�V�I�?g�f���\X�<����8��U��Ĭ���^W��C�G�p��h}Nw���}p$_~R��Υ�d[g���+�J���q���U��x�6�u�XX�M�Nv�!�`�(i3зq8�Ј'���Xw���,D�������D��u�(n�����J�q���U��@����gG=%� g�VvO����&{��X�/R�ό���.�}�
�?���)�δ��Iћ<���n`5�fK���ġC��װ�:�iԟ��=��.wd���/�t-gx��P�\�<��R=p���W�.�Ӂv�u�o�\�rG�,r�.!�`�(i3jݭ�F���X+�f�f�!�O��1���Sns&���)�δ��}�\���;�YǯXan�M�:�����L5ӥ���98�
x�?���~46��E����FkѶ���� �G��:�lL��:�iԟ��=��.�{�s�*���%�T�t��{�G��ͫ������:[�F��#������+�J��;�?�կH��%�T�t��{�G��ͫ������:[ۚܖ��`��AW˟����V�����lJ��I��p��mK�������T�-07���wұo�35D8�y�\6?7���6��v�����:(�B��N�f��-yMc|Q�Xn�	�%��6�S�C���m���d�hY�%Ͻ��Xy|�W��$����>&S�XQ������;�oz�� u]�MPŪ�\���S)����LB�g�RMm�o����\=u�(R\֎u�D��u�(n��K�f�1���~!�`�(i3!�`�(i3��=�$��mp�E����!�qg�XJc���!��{*9����*��� �iK�D�b=����LB�g�RMm�o����\=u��\���S)��p�:�F!��D�����k$ !�`�(i3!�`�(i3٪�o�_&�&H�y�66M�Z�i���&|�N/�C|0���f1�.��N��X/�7�{x��O>�7�,��n6�o8:4�I���c�90Mj�dL�{y����i�q,?5qr4�Ў���<�e��BF�U���e��d9=���u��r��J���hB;PB����A����;q�"��ӌ�r���̰�!�Xy|�W�(�[�*n��뾦��#�-�p���p�:�!�`�(i3� ��U�_:��}Dq�f�o;�Ul�|�Ƀ�?PAn�#�7�;�j)����r^*qA����6\�4�@�� �-j�1tSjv��o�t��D��u�(n�D5���.p�YD<=���+���q�����̰�!�Xy|�W�(�[�*�ۢ	:j���k¶lW�x��7��PB����A!�`�(i3��X�zl�rx��E�x��7�� �����2�w����6��j��8Tʈ�Ym�����xb}�	76�&�� Ӗ�t$�)�vx4����!��:W̘
�6��j���