��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�-Q3�Y-ǋ 4�i� ������[���a�8%`��4�s�6�XAoeuxLZ�#8������^F��W��`��9����`,��I�|��]P*m����)O��Ξ4�"�\�� ���K�O�{�����8�\�3��>M[c\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|����(Ҝ��;�0��'>=���uH�!���Ȗ��h�}�{Sh0�.�	�Z���}fTV����~�hbHp|�P,N��!�Ψ�	�ǳ۱��@�QU3(�R��W�ew2�\�����	x]̍��;����?��|:�-gc�n O�HߵgB�T�V7���p^#����*
��$tU�U>r�O��C��0��ד�̟a�,��I�zb�Z>8��������]�\������������;�kv޶Gl�!��TN0N��\�4�si�W���Y��݅ 0�1���جچB�)oo@���q�&p�`�������N4�$�����(
� �AH�T�t��3��e��ME
^����c�:���0�F@�4%�u�L�r��3�jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��dI�ZS"J��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�ĲW��,)i/-�#�v-~x��䂁!�o��c��(r���U��� ���yX����!���b���q���1�:�Ω�S�T�;Ϗk[�^��_���ˊ&;�@���,������0�=j��S
��.�z,y1}Kط��4q�������o)�]rR��ӟ-���r�1���X���`��Fb��҆7���ө�q�#���Z�>)��<H�-��*����Kp&�@���k���a�\����9�	��%ι��QG�����U��зq8�Ј)w�<�_N���i��I<��fҾ��9�Ǧq��G8��=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A�����
�����Yl���#�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��kv޶Glbq�Z��T�I��w��,c�A�L'Qī�*pY��?� Zh�RG�p�PR��{�&�8���/�2�ZwŃ�9��|�����|g�Y�'���Xwp����B<�D-Ε�(�
t�ژq���U����?�"�,�>E����-��%Mό���.���|��p�}J�A��j��\w��0]%��C���]M��_�\"e.��xu	�*�QN����q�1Ig�I�?g�f�P���.�V�k�J'�����N<���d�k��Yu>�G Oag�qod�֓��+��T�����TS%�}< V��Ҝ��a�N�}��t_���Յ;��n�a�x�a(􆿳��Ak�y�y/��=��K��]z�Sk����+��_�F�����CY���<�;�L���9��Xv7�je*���W@�$C�~x���yM�y/u�!]D	e*���W@A�;�֋`N��7�j2�٭?(Ů�C�*ȉ�Mx"��������c�A�L'��!�a��5�%]���a(􆿳���2����.���N����]�u+J���r�S�ML��ʐ��$�J��u�v(Ȑ���,��P"G�wk�١��	;q��^̽1��R��ӟ-�F`���G���`y����@����gG�?#dK1"Sr��3�9s&uA��f���,(���B��ɓ�~Ҡ	u{ᵿ�����"X��[��Q[R�7}ϼ 8�����z���	F��6�q��T�ٮ|�,
����$C�~x���yM��?IK��y�8���/����,D$ů6j�e���;q��4��7���b�Bϱ���w�K�})9ͬ果�k�V\���"X��[�d�a�4$�b!��u�^�9.�JQxZ��j�
�iB{�Z�_��?� Zh�RG�p�PWȹB:�Y�b:m�X`�7���ө5�_)��A���`y����@����gGT���/ �c%ij��d���0y�	�C�u)�6�3A�)Oq87{�Z�p(���B���ި���������f�T�\ ������q�f@z���Q����\��2��� L�>\w��0]b!��u�#��?@�]зq8�Ј'���Xw���,D�.���h��Sd�[��d�٣���zR�K��I��� (�\Xɵ�y��`2����]'\gWg��	�Z�kfc�?)zni��`���φ��<�6��jf&�~�7�W8�C���'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g�'��o�x�S�ӄz4/s�1��p��nF���<�W�.�P�	��
�Q�}��=m緒Sr��3lr�{��|e��0�U+�qbp@�,\ͨ܉p�T�8���ᛚ�z�Ji���nF���<�W�.�P�	��
�Q�}rI�F����ez8�US�/ ���we��0�U+�qbp@��x��'�^_��Sz�t�!�`�(i3%��v�ڹ߆�p�h��d��JXl'�T��~��?u��C@!�`�(i3.�
9� ���(ٗ.;���JTv�䵶
�t��T&��ۥ`�M?��y�!�`�(i3��_	��Eʨ�`N/�J�J�~>EX!�`�(i3�c��;C �3<M!�`�(i3@�c�*j2⎜ä� |��&-���xԾ�J��RQH�RtV�^,\ͨ܉p�T�8����_����,�d��z���	�/����*Q!�`�(i3�����!�`�(i3f���8�67�|g�)��E�g�������(ӈ���m�r����
�:qEp:䩒=]'!�`�(i3@�c�*j2⎜�m8�� &-���xԾ�J��RQH�RtV�^;�jmT�#�#}�{��7�i'����^b�~R��ӟ-���J��RQH�RtV�^!�`�(i3�kv޶Gl7�|g�)���h�G KH�����j�/����*Q!�`�(i3�	��x��ݚ�Н��B�'��a�
�oz˸�1�"�����nF���<�W�.�P�	��
�Q�}!�`�(i3�5ߧE4��!�`�(i3��Ě���ž_�FȮ� л���S�	RN&*�8#u���;�jmT�#�#}�{�@�m�W#����p&1"G�p�P�m������� h�ҩΟB�'��a���p��b���ez8�US��h�G KH�F;p�	p�r~�h��ݚ�Н���w�w:�!�`�(i3hs�����F;p�	��Bf����{_8�Y��=�}�Vݨ��}Dq�f�HN��R��F F�E̠����l��2l��*��Sr��3	-�L��&P��7�j2��S]�_�_��u��r��!�`�(i3'-Bd8il�e���;�̓������x.�Knq/�r�]/2�ݚ�Н��q�9�ͭ�M���V����Bf����@h G0L�[���_>������
�:qEp'{w#/ B!�`�(i3rI�F����ez8�US�E�g�������(ӈ���m�r����!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�<�6�Q=�x���y�d9JR�tŸ3y����s%lPb]�g��X�a!�`�(i3\���;����j� ^�Ks!��f^�j)�UK�ƘpK�9�b�T�8������R��y�%�j��LaZ�?�u��r��!�`�(i3CTm�q3��;���b�t�d�l�K!�`�(i3�5ߧE4���ݚ�Н����F��O�VA�ڦ�c4�5ߧE4��}�	76�&�j���Gp��ܐ�}�)-��^8 ����j6ۮ�m_	Q������m�͑Q��8���
�oz˸�1�"������c(��BԆ^����ȕq��N��%��T%X�;3�#��j��Qv^��F;p�	�j�q�7ר ʋ�a�Jw��3�Jz��X.	1S�#@F]'\gWg��~ޥj�!W�.��|ȃ��!�M��9�a>*<UB3 �~k�%�������&G�H����o�γ�ha��o���zM#��m��k��M��� ߌ���*`2d�爔�C.�u�X��I�ՠ���7D!��6�G�CQ�}����l��M��/,;�.��1���-����!�`�(i3�L�s;SF`R�"�ѧ!�`�(i36�&��=�K�o���,X�FU9Pi޼WaU���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��8�8!s�����4��;��R.���U��)���Y;e�iKI/B޾Pb�i0[���S�J\7CZ�zk��X��%2�/�C�7�癆cgQw�c4~Nr_�mS8<�n!�`�(i3!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"�[�	���8���N�C)P<�ܓ�YE�9�ؕ�^3rdS���q9+t�}��=����t��p��b��!���?t��my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�$XR�QܛOcOZail������&G�B�'��a���p��b��,�NQ��.Y�{'%s��jb�ܳ���p��b���ez8�US��:5A��p|D
�W�ɪ
�oz˸�1�"���*8j��4	���_�239@��C2K���l��#��I�XƤ5_���Q����ݗAn�W��B� �b��!�`�(i3�>�u��8�m�Qrx����NM���fĉ>99��A0ok���H���������A�}p���I
�����&G!�`�(i3���N4��?���_e�� 0�.3�!�`�(i3�5ߧE4��!�`�(i3�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��pɒu��T^�h\�%(㷾�!N�'�y�G