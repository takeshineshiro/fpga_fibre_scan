��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� (� ��"fف�������J��.���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:����>�ፑ���ԛF��W��`��q�©��7��#!l'���h�W��!��CR��=���u��N�w	*D���y&�f��+K��[y��ڂ�Vs>�+��T�,F���J�/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&���7�os!w����]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�K�MV}xj\�iW�(� 0�D�A~����p��ؚ�fD�~����pn��-�4ڭ	���
��M!�nz��m��+�ڔ�wV��y�p�cP �����-ǋ 4�i� ���������	x]̢/����w�c.$���S���bJ���<����PГ����"��N�� <9[�8@������G�٘���ty.hSN�����\�4�smg�:�TZz�0Q�����F���0FUR�.�;�~�MUs �P�^,�Q����j�_��l�؊9��8���M�3)ͰnL
�k�8���҆�|n������}�K-���W}��@_���J�Й�m����u�����w`q�tc�ؑ��g�=Iĩ�m��d�7�Q����.P2:}��>�,�_'�hQr�k@Q��j��C�뫰v]uR����Pl����N�Er��xXc)O�%���ʅ�$n��RL�a)�ƞ��U<���G�/9Ɗ���ބ�F=��?�r�7C��H���j�v�?��$m��2߼
�d�
 O4�J�|(�����	x]�<���eo�l$����Pfg��w{��������PГ��-�������n�GE^��.�Ū�'E���f!ۤՀ/Q9*سBK-����s~�j1���u��w)�S �J���vy�~篟|�<8�F�-:�0��E_}�8�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A�f��Wj��y�͌�4r�O��C��0��t�z���� 0��]��=��c��v�u���;�=�I���ĭ�D��)/�F�5�_2��VU(��z�j�@ȶ�h�..��X���#�}Hy����͙3����w9J��[g�������t�5O.h/�o����Rw�@��V��=�L��ޖl �f6�u�+��e4,��͞N	��;�W_)O����d١�����m�Sb��RL�a)=�y�~ N	:.���nX$j&a�"�A'�_.�TZ�7C��H�y�ƴA���e1��=q����\�_�?h-�}4���Qt�j�1w>�w���������U��֊���}�cz�m�!=�y����h�}�BK9�H�.�c�T'9~�I�Mc�o?�M��;]�u*z�f��U�0�v:�MS�i�>b�8�e�
uC��%�e� �0��}��0w�\���J�����\�4�s��Иk@D�Bg�3���M Ce=6�([6�?�W����7C��Hwɶ R�p��4�s4�o�qR��p������M<D�7�s)	w�N\`�a���!4d���-sk �0%̄sb�� bL�k>F�泂�0�V�@���RL�a)zAY����-c�J�M=�2��&�m.([�G	{8�:r&@�G	���su�]bu̎x4�J��|���>�
� �AH��>�H֞ T�{ ��ʥ
���A�8���Rk!1J�Й�m��b�)�� �G�q�����-���p/D#r�O��C��0���^S�kUC��._�U�����gP���)�$�ɀ�&}Xa��=}���mb�.G���6FO��fҶ���S�X��Z�Ʒa���uSz�ޚ�����RL�a)��F>x��F���f���euw���wB"l��u���;��I�6r��f-Ӵv����N�Er��xXc)O�%�!�&��{G�3�^7����$������@���F���<r�O��C��0����bm���?��~S� �.*�1=\5�"3��
f�6{�I"UTG�{6�m��2�ӭ�D��)/�F�5�0`��E�%Ct�Zi���u��w)�S����w7��Mv�9NFgӦԙ�$����џ�_�v%��ˠ{�t!�.�r�c^�e���zǒBs�&���b
� �AH�W���,2w���$�cUY��p�5NJ��f���F@�4%��]��N�"�<�/���;c n�b
� �AH� K�`A���vJ�^ <.���f������$�J�Й�m����
|H?S⏸[��[{��$')Y�8}�r�O��C��0���/���k���_0'Z�Q�%	�u���;�4����l�~���&�����d����OX�5���\�4�sR���i1�TT	q��$듍�E��WWSt!K� �~�MUs �ˠ{�t!�.�r�c^�e���zǒBs�&���b
� �AH�}��� ��� �b5z�U�՝!h�.���cr7�F@�4%��%dZ&��Ǯ"�lf�~��m���w>�K�6���	x]́��D񛎣��]ewk��y�'�J���<��³6�&N/���wx
d5�(7���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�YZY0@ìO��3g�ݜ��s8[Z�`
5��*�zM�D_���.���nEA�i�+���/?�s�m/C�N{a�9O��Yk"1/a��ʁކ�+��T��٤�2[51g���i��T!ea�8���A��>s>;�.�z,y��}����E���ƪϤ�Yk"1/Y#_Wӆ�q�©���H��JnXeS5H�j.F�YZY0@ìO��6�g�m��+5z�P�_XV�>!�/�7��u���nEA�i�+���/?�s�m/C�H*�m��/2�ޅ���?�y��h��ؒ3����]ͧF���y: ��˘磋��w.V&��B֥�(����5��-��ˋV�{�j~�|�ߦ:`�'ࢯ9&xc闑^����S����ީ��ƭ�����'c��2�Ặ��Ϊ���Jjz�^�R@Κ�2���ei�b9����r*�^�	�����\{F˯�+)���u*K6HT�����N�~ `�T�v��1���;ε��IÙ=�H<z,Ҽ&�jV�{+穴ʐx�?�'n�^0o)�X��2S-v��B��q�T��&�����-N���\�v�T?�7G|`^�R@Κ�2I��RhF�����<ɣ�'n�^0o��~+�ݗ�p�ϵ�DE�~j��[7�d|���XP���)٠����g()��ikp���H����[7�d|���XP����@PVڵ��#���F<�r�5j�'n�^0o`�U+�PA�p�ϵ�DEG�p�P�� nU�IÙ=�HF���m¡h�5,Wl�/�O'�=��� nU�IÙ=�HF���m¡h�5,Wluϛ�?ud�[7�d|���XP����ŗ������U���gFck
���/d�s��p��'n�^0o���˟y>���c��d�|ݔ�3�(n�'��b9���:&�>��s,Y�o�a�gf{}#k��Ȁ`�>:8�A�/�����%>%��"����?e��G�K$x/��&���7�ܥ��2�]Hf��?)���v���H�息��yN4&��M	�D�$��띂ii�4];ˍH��T�K"
�Q�͹�Ɩ,���#>c�b��v݋N������M}Ĭ����[7�d|���XP���Ý��'��fÁ��/��F��H��\�v��_�R�GI�~�џ�.���hGD@�F��q���i�����Y�V&��A��.D�.���hGD@�F��q���i�����Y�V�~G������"�4];ˍH�:(�������҉�}�g��iW����<5�;������*8�4];ˍH�F�� g��³��wQ�q�o'�4];ˍH���������ERF�G{؍��R��j�.(Wx*��|��pe���b�c��Et��q���U����?�!�`�(i3��|g�Y�'���Xw�E�i�m}6	��	Mk�rv�ј�"��Z鎬����A��:6])�/g\�H)��,vw+�ne.��xu	���S8����ٺ?��Ʃ��6��G"ڻ^!�g��U-�ee�@Rv����my$�N��o�/���;�%ؙ,{F�"�,�>E���TD��ό���.ӈ�=�$��zigzA=v)��(�
t�ژq���U��ꢤ�OgB�Y���c��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<�(�&�q���v�ј�"��Z鎬����Ĺ#{���4��}�<������K�]2�y�Z鎬�������(����U6�bL��W��_�ړ8���/�����FZ^�u:��_x�����	Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/�I<��f��tN2s���(����5��-��ˋV�{�j~�|�ߦ:`�'ࢯ�Ah$��>���67�a��c���}��D���(��z�j�)�q��1�:�Ω�[@�qR�� (� ��"fف������G�p��0��L�r:Pip<ɯ�nv��2������開k����6U٤!Q
���g��Vܙ��t�cُ�Ջ6�x�p�=����w`q��La��Y�E����m�s�*�MOL�ӯ.���w7G�����]\{���bq'���7�-���+&hJ-.�{�ނw�?�b�>޼�\�vŕ�`UNP� ��b�FP&�5�+�zL͊�q���0EQ�W7��`���߼
�dgn�*�Q3#*�ۍc(y����>�g�R�@�6�֐����o��TT7���1���P��(*� ���Y�8 )�\�~xy�֍z����I��'�3bQ=�3��� �?́Ặ��Ϊ���Jjz�p�m~|����@��T
��;1z�}�=Ll�����,۽���dט�w��饋����Αǜh��6���C	)�H���o��qo�:���$��Xo��yذ��tp~z�r,Ln��S�W� X�6�]\{���bq'���7���T;ZJ5�$��Xo��Ȃ�u�.�1�a-���7a
��r�Ln��S�W#w���	(���B����_T���a�aq��hx��t�#���F���U���(���B���Q��ǺΕR��ӟ-�� >��Ȼp�m~|����� �ܰ�a\Y����)���8҉g�kG�#JHn��z������W/S��8(�E���Kt��嘦"?k��g�,P�n�|��{�ru�?�=�r�@^7&ģM�'n�^0o�<:�W�_�l�J;�Rg��dT�W/S��8(�E���Kt����ӯIJ ��`y�����g�,P�n�|��{�r1��j��Mشˇ&�,�>п�p=	�˳͠m�xW��9u$d9��}ϔ��J�s���
�k��!a�tc�&ck��};l�-���L;Л��|#9���hY����r�;*�}Ւ�~ܔp�l
d�o�R�N:��,��g�7�s<��MR�������c�A�L'��!�a��5�%]���a(􆿳��?ƾ�؀qjZ��H@H�֦g�㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���o���ia���lC��U�T�\ ��Z��| �Ɛ�5����`Kw¹��<d���	fdLn��S�W�כJϾ�i�I7��-5�[NESeV�q8M�_�4�|*uN�wHZr��AR1<�N�؆�B��W+`�x�oP��@t�&�e�5
��Ib����rs�i�jf� l�Ǜ�����e���%ޘ�g��U-�e�T�'��k�5����`Ke,fi�U�ž�'�t_�GZEh5���'n�^0o�hŁw:����v�8:��|`��'J�	�LÆ�c�9ʼ��$�G�nJ `1	�<�����!�F<�+P���I��ž�'�t_�B�uʡ p�m~|��;~7����WF�r�f�t+Yi=��o�IÙ=�H��w�K��b�����(`��ү/�O'�=�eX�
\;�M +�gf���a\Y���c_����+#��.X���*"v%)��Qcm hP"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y���p��nk�r��VYW\y]/�qF+Yi=��o�IÙ=�Hw¹��<d���	fd��Q�b��3R�^Ƒ���P4ǲ p\匔'������^[_�e��IÙ=�H��M���o�G�m�?E+���7�$��Xo�e_�d
���ݪ��1#��Z�����XP��ȗd�uY��K��T��p��`�Q;?�͆�%l9�e\EV	�*�����I��'�����Dɵ�p�AJ�e�$�^[_�e��IÙ=�H�S��?��L	�<���BS��nH�W�J�S�̧���� ���U�e�7����	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�����NlU����z~���ӯIJ ��`y���p��nk����eR�ʨ��_�\G�k�y'��aLn��S�W#w���	(���B���Q��ǺΕR'),��`�LR�Ssnň����T%wxE���8�V����8��?�d���&��뷖iU�p�m~|����U0����d5�:�w�+���LQ��b9�����:�{��ߘ�)�I�3�"��+W���F�^��NPC=2崝�Q�gL#A=�����ׄ�+Yi=��o�IÙ=�H�z~~�Y_" �g8Yw�
��vK���w�K�b��2W hbvk~�#x�%��4�w�$��Xo����BɊ�y4<��!I�Ki0j@$��U� ���_}U���x�.N�DMY����U��t��ܣ^\t�*�00?�9�f�u:�]X��w�3Ɇ��C��ǟ0�]ov��Kԟ��j�釸�{�~��U�zGСi��ޕ!�\����[��g�H}Ct�U�)YB��|�L*.>�+S�+8@��31U�Y��-�E#�墙������6yT��GY�<7|'6��}������lD���7|�W�q���Ì?���/�\��5����`K��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#x�l7�l�r�#���FN��H4�[�S��'������bpQl��u�!�`�(i3"�,�>E���]�!����w�Հ��Ed��>�^���n���g!�`�(i3зq8�Ј'���Xw�j�7����`�z��Y��),�B۸��L� s�j8����DzL��k]m���޿�*rM�W���D��g�[�$��X�՚��l��Hr�<Uee�N�����H�OM��`�@����gGW�RJ����@{2귑��r��f~T�􇃬Tk`�|��K�z��@d��שI4��欱���j���-+��B�G�
�CӞD���:�#�.��N�x%�%�T@�zF.ZVRѿUJC���d��ݷ���r�$����v�b!��u�9*�"FP��� �mD�eJ2@����c�SD�=So�?D����y(�\��`8�(6�@����gG���:��,��!iJ��?��(��I@1���t$I+��f�kN�ı*�7`����\Z��K���BE�B�M��GKY��B2W��4�`#�̅�\ ����DzL�#�r��8��y��?{�%�*ܑe�W����n�4�`t��D����M����A�m�([}�@��L}�
�?��V5VM�d��LX�Y�k�:A�	S�r��AR1<��J�@Ym��`�z��Y��),�B۸��x|qj0�vے�(�iF��׿]�/�˟��7<���������	N^�U{xN��i>r�<Uee��~j��6"���T�@����gGKCYb,�q@9
!�gwe�ŉm�m�jp=�>��o�
�v�ξ���Ix���KaIW��d��ct�:��RE�QS����>��"X��[��Q[R�75�e`��9��əS\�
���X��d�٣���������ݹ�0���f�Nd+l�Yҽ֗�)�|����P�%.^F�	��lC��U�T�\ ��i3�|)sՀ�23
����X%�(�ƇBHx\�'���Xw s4S�'�i��`�z��Y��)h��{��Ē̫� �[:�������CyW�f�tR�wX��J�W��7/ĩ1r����j�1зq8�Ј'���Xw�j�7��ct�:��RE�QS����>��"X��[��Q[R�7�
�CӞD��m�q�/�Wv�A���d�٣���N N�S��M#��W�}�IUr��ӣJ��
�|D�of�7���A3�(N��㎏qló��@d��ץr�&U������G|M��i�ܰAb!��u�R���V��"���q���/y��g�'b�t	�U���C��O]r�<Uee���R�}vJ^����`a�ct�:��RE�QS����>��"X��[�d�a�4$�b!��u��Ɔ �����Vd�+k&v�IzZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕?��`���in���㬺ƃ
ᾆ�x�T�\ ��i3�|)sՀ�Oi9L�:�k]m��KгoHG�K[�x�X���z��N��ξ���e�J�Pn\�pD��ZOUi3�|)sՀ�Oi9L�:,�۞��	���/y��g�'b�t	�U���C��O]r�<Uee���R�}vJ^����`a��כ��p���lC��U�T�\ ��i3�|)sՀ�Oi9L�:�Òҷ^�vW���D��g����H���	N^�U{xN��i>r�<Uee���R�}vJ^�k��76��&́�������n9��g�剭MaG�@y�a�P�Fpwe�2l��4��a��se�ξ����l~�U�n��(���i3�|)sՀ2��2,͕�%�]�
ƇBHx\�'���Xw s4S�'�i��`�z6/��������рӚx�Fh6�����ݪ��°������R�wX��J�W��7/���_�Ps޴�ik]�7A��(�n��rs�i�� ��*b�+W���F�^�Y�7#�xI��;mQ��8���/�I����"�A<�}	����B�[���d�٣��c�A�L'J����l�!�+���LQ���"X��[��Q[R�7�n~�x��<�,���E���Q]� _ό���.�}�
�?�)HVi�pL�+�@'''���XwI����"�]^U�*�!�$�����P"G�wk�١��	;q�U���3
�v�v-}�	mp����"���;���N~�y��l�6�T�\ ��i3�|)sՀ]^U�*�!�8p�u�dS�P"G�wk�١��	;qJX�D�0a(􆿳���2����.�ɷ���/s�1��pq��T�ٮ|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/����,D�;��[TM��s�hd0AԢ�a\��F�dH�Dj���G�Օ��qvdЧ^{�j����#oM|#9���b!��u��d�@���Gғ�vq�\[$Q��
�̞��>�nQ�rV�}!�@�?0a(􆿳���2����._�i�c�/s�1��pq��T�ٮ|�,
���Ϊ�/-T)x�?{���x.�Knq�z���a�R�wX�ո@����gGWm?"<���Z�n�f��Z鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀ�T:���V��%�	2��d�٣��c�A�L'J����l�!�+���LQ�M/^���iq�VD�Lg�q��Dv;g��"X��[��Q[R�7�n~�x��>c��?���Q]� _ό���.�}�
�?�2VP��Ѣ���t�Yǝ�b�Bϱ��ᵉ3��鑘2����.+w�7�
�p�	%6�n`5�fK�\w��0]b!��u�����P���+�J���q���U��@����gG������0g�z�&��Z鎬������_�,�;�7���c�	4��t�f�d�٣���N N�S�qg2�K?\�E��ȷ���n`5�fK�\w��0]b!��uፍkv޶Gl%,�6��Y�]�!��	Ǹ�y85���ǳ@�M�H�ɇM��lC��U�T�\ ������q�f@�]�gv���J�����d�?�V�^�E����FAԢ�a\��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_�k]m��Z�����h��lJ��튝�b�Bϱ���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X�v1a{J����%]+aúAV�!s���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�G9�:Q��Ĵ��ޯi�-Qq��PnO�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv��G7```+�!�`�(i3�E����FAԢ�a\�y�T�g}�Ӄ�Q[R�7�����bpFn�H�~M�!�`�(i3!�`�(i3xZ��j�
�iB{�Z�_��׉p'*EF���L��b��v݋N������W)j��T�\ ��i3�|)sՀ*�şxˏ1��o\�B/M����*�зq8�Ј\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?�K�\7}�W, D�cg�}�+G�}�	��U,�(�)8���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�[��m�U����L�F!�`�(i3q��T��J�s���
�k��!a�tc�&ck��°������R�wX��}�
�?�K�\7}�W,��+G��ܐƇ:Vxp�k�XLF�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.�>��왩��k]m���E��Y��{Z�0@gĐa�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D����y�[�%��g:���
A�%�q���\� 8�����0y�	��sC宸I))����A�m�(/!���La����-U �ZJ�hEc�>T3�$�Y��g��ZR����z�Ji����^.�]�|�,
���N������2(wUF�|��: ��ao.\C�k��~��Kؓ8���/��%G��ly��!iW=�!�`�(i3!�`�(i3�E����F�ANʂ�g��U-�e^��hדܳ\����%�Cj�|�{'�v1a{J�&��	�>��E����FAԢ�a\�D�����R�`�|��K�z���k��$a(􆿳�ټ*w2�56�����bp�WdM4@�k̇���A�D#�"sO�=�ͦ�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.�>��왩��k]m���E��Y�"����5�Wȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g���j�|�{'�v1a{J��9H�P�.�"�,�>E��P"G�wk��r)��ׁ�a\Y����)���8˩��F�{a(􆿳���2����.�>��왩��k]m���E��Y��vc��W�xZ��j�
�&�j��1�a-���7a
��r����~v����"X��[�d�a�4$�b!��u����M���X"�,�>E��P"G�wk�١��	;qBvGޣkQ�A���ۖ�k�V\���"X��[��Q[R�7d�x� �q兄�`�&~�E����FAԢ�a\�/��A����Q[R�7d�x� �q���
y���E����FAԢ�a\蟱�c��qVwRD§B ���`y����@����gGT���/ �Ve��˅�O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����Ed��>�^�����-VLy��Fp����L�de��-@��F~*7���&�_ƃ
ᾆ�x�T�\ ������q�f@�]�gv���J�������ߧj@Q�������f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/����,D��ǉã1X�v1a{J�Bz��s�V��8�P��Ά���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?��I�_Pg<�4���TS3��v(�y�xZ��j�
�iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��Q[R�7�)�`E5�j�W�����ד*(�]F�5���V���F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����]�gv���J����0;�����q�:�"��f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/����,D��ǉã1X�v1a{J���Ꭓ�[��Wxu�VZϫ��0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?����D)��ʱ�O���E�`JcUȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����Ed��>�^�v1a{J��vc��W�y��Fp����L�de��-@��F~*7���&�_���/���l���F�8���/����,D,Q�\C�/�����C�V���3��U,�(�)8���0y�	��sC宸I))����A�m�(};l�-��'������݃�Q[R�7�
�CӞD��m�q�/��v1a{J� H~�ɐa�x���w�K��r�]�4�P�l��=5;R�ˊ	18)Dg�|4��`y����@����gG,#�g��C�x!�H�Z���,�q��T��J�s���
�k��!a�tc�&ck��};l�-���L;Л�����Øf}�
�?�N��	�Ȓ�cЉ�M�G,�A@�Q�y�� Y{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Be��`M��
AԢ�a\蟖�S� ?�0��E|�,°������R�wX�ո@����gGQ��6��'�iA'R�	z�#,gB��Pߺ0��A���ۖ�.Q�2�>�f���,(���B����: ��ao.\C�kHgN�����`y����@����gGQ��6��'��o\�B/u�:o+���	�����aq���皒nb�B�f���,(���B����: ��ao.\C�kHgN�����`y���h}Nw����ǉã1X�����m�(��k8!�`�(i3!�`�(i3!�`�(i3!�`�(i3�k�XLF�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'؁C�*&#�4?�o�5�h�B��A�	���\!�`�(i3!�`�(i3зq8�Ј\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?��x�������E��0�Z�7W�:��G�z㤧{��z;#o"�I0���ԏc�r�(���ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_�E��Y��Q�
w�8F��6�!�`�(i3!�`�(i3!�`�(i3���^.�]�|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[��H	X��E����F�f���,(���B����: ��ao.\C�kHgN�����`y����@����gG����<��y�@�v�&Sq�a��z#׊;w!�`�(i3!�`�(i3!�`�(i3O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv��JeYSWe^E˔ �y=k�2�u���e�՝*U�޸I))����A�m�(úAV�!s���0y�	��sC宸I))����A�m�(/!���La���Øf}�
�?�rS������A�8��|VO�⅘��a�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X�v1a{J����nFy� �_Y��t��3
�v�v-}�	mp���aM�v�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.JL���Z'#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#x���Z�"���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?��I�_Pg<�(y�.
جH��O��U
hPߺ0��A���ۖJF���@��a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀCeFJ5x�_�k]m����DބiM�YG5`FFB5=��)Q�ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g��սÕB\�6N �S���}�cЉ�M�+!�j�8�3
�v�v-}�	mp`g�_��iB{�Z�_�1�����\�H��/Sg޶��j�}a�cf�g��U-�ez�r�6JL���Z'm&����T��Ŗծ��7W�:��Z���⿳�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�*��/qRr!�`�(i3!�`�(i3!�`�(i3�@����gGQ��6��'�G����1�E�AvY�5�h�B�΅o��~v��a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ���sC���X!�`�(i3>�3x̪�1�]�gv���{V�-_8���G�7W�:��G�z㤧{�E2p��F4F�[��
5���١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.JL���Z'�ɴU�ԉg��h�=m�(��k8зq8�Ј\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y���!�`�(i3!�`�(i3>�3x̪�1�]�gv��L_v,<=��}�I����&Sq�aQ�y�QF��fK�Ěk.ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e���B�/J�W��7/�CeFJ5x�_��DބiML�瞩w�j���@ΙN�)ɣ'�ikȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e���B�/!�`�(i3aZ��qA�E��ǉã1XBz��s�V�r�G� Y� {l��	�g�yl��6��������hˉn犫��0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX������n�I��'��Z�<��H��h �=�%Ah�%4
>��XP���ϝ*�yo�2������}���z�78���it	�Tߦ^Cg��)1�q�ܲ�xΠ��yGb�X~�$�	�hbvk~�#xnůc��o@h�5,Wlr�r%)cA�-��h�m ӫ/��m��?�4D+w�����������f�l��=5;���wGu�ܝ�s2����˨(�V�֪��o�� �}��2m���l������L��@X�hD��$_s����z2�v�~�g��27�*Y=���į�4 _;��i�1@�f=H5H�n��cM�r�z�IF�@����gG�XpAS"Y�j�`M"�,�>E��P"G�wk�١��	;q�� ��-�BM�ܤm|�8ɂ�T�T�\ ��i3�|)sՀ;�7���c�����-ќv���z�Ji�q��T�ٮ|�,
���A�;�֋`NY~�y������̡99��: ��ao.\C�k��2�l��
��"X��[��Q[R�7He�-�c��Y���D��3��b�U�,�6���'K������V5VM�d�/|�;{$�WaU�����W�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �2(�����N��j�'�c��?F�*���#h�3".t�|6
�Ԟ-zq�^�W�	mɋ����Q��ǺΕ�A�m�(F &_{ _��s�֙4�(�Ҁч��>�{��u�Y�KG�[k�|�G ��Y��)h��{�����R(�.ָ�d���!i�� л��2V��y{�~7�S,���n��_���V]}�����j�ݣ�heQ��O�6���?l��fN���)$���R'+�^���VA�ڦ�c4K��l���V��J��n������~��_T���a�aq���)�F��Օ��qvdЧ^{�j�k��L�ظ�d���!iV�Ո��+5�4��c�.����^_!�`�(i3!�`�(i3G�<�v�W�t�3���2{��	�!�`�(i3ϟ��7�4Ï�6]S*�N�ǁ�f�TpD��ZOUg�w�9���+5�4��c�H�v�m��Y��),�B۸�b��?�GޮHN��R��?�d���&�^�a���3�m�G�]=t�G��!�H��n	l�ۅ��$���D��8�tufJ*�Rs�08�b(����X�zgz�'�̗��������p����Se���7�}�!��P� d�c�m�/N0
��=��9�&g�{w���z�+��@-�-'͏��������X�%?gV��U�x�l��1:�N�*�x!�`�(i3�
�I�>y!�`�(i3���u�UgF˯�+)��&�C�/�zg��p�r�X�<\�!�`�(i3�{�BaD�A���ۖ$����h�5,Wlr�r%)cA������]!�`�(i3��'abW�5�}�]���rQ�4��+�]�U��y!�`�(i3�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��� л����K֫ ��")�/K��sb��ȇV��[g��z���.��!�`�(i3WPtA��ro��� zv�۲=�k2!�`�(i3gh�䊉�䞘gx�n�W�����v����?�e����kn4@Q�/�!�`�(i3�_F�k-��苇��Fe#OOJd֯!�`�(i3���ꀍ�˺�Q���f�?ǉ�=���%>�rG��M����{����"!�`�(i3 �@��&}��{��W�#�r��8��n咫���!�`�(i3{k�h�+d�/Y�Z-u�}#�U��X#�v�%2��ݚ�Н�c@��;���ז��6_���������I��2m��+�Z����y��3�z?Z�!�`�(i3�,\ަ�It��+g[�!�`�(i3����$G⃍�����u~xgA���������6%�a!�`�(i3�gCu(o?C!�`�(i3O(�i&�Q�J*�Rs�08�b(���,�7�%�aR��ӟ-��1��NhO5!�`�(i3ΡKCh��(	�G��^����K�7��I6&�H@��!�`�(i3$��:�e�hfH'��!�i����VZDf�?ǉ�=<�6�Q=�S�'���� ����}`�/��+�!����/wފ����!�`�(i3Ta�F�O���^�#��\�'�ݚ�Н��K�^����\_9ͫ��Q������(���^�,\ͨ܉p����O,8�ݚ�Н�3Lv	̅���X;p`�(�����!�`�(i3Gظ0����t�%�Z?��<�ry^�
�:qEp��:��Zg�Hn7�(�!�`�(i3[�л���7��+��΢t�3����%�toqP�N�ǁ�f�T�A(夽�	XT�1!�`�(i3p�n���:��]]t�GR�D^f�Nd+l�Yҽ֗�-T�"�N�ž_�F�w�R���y>��yС�[�(r"(VA�ڦ�c4��L���B�@o��[ea�8��������?9|[�,HJ
a�\7�"
q����Lt�iZ]XF�hx��G��!�`�(i3 k��v(�Âv����Y���a\Y����+���LQ�f�?ǉ�=�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=j:�Mpp�}�(�-lc4�j
Թf�?ǉ�=��X�u��
)\Y����4MT2g�ȨQ�?�Q!�`�(i3���ȍry��	SƏw0��П�+�
8'���Xw�j�7��9*�"FP>����qZo����!�`�(i3/8«E�A�J�e�!�c�A�L'D�g�=a�iA'R�	_yZ�'lN$VA�ڦ�c4q�\E��0�aR�J�}#�U����5�W@!�`�(i3�.C��ar�=k�Hg�]T�o8�ժ*)xJe�2��}��M�p}��ϟ��7�4�Mzu�P�v	��Yu(�������e�-3���9Q�����ݚ�Н�Y��
�iC>N0Θ��ݚ�Н���0�&�ͭt�%�Z?��<�ry^��������c����҅���H5t6F�7���lJ����I�?g�f��Qө}�_g�?�H���w�1%`Y��V)�%?gV��U�x�l��1:�N�*�x��'T���+�htO!��nT�Ā���-@��F~*7���&�_j;��q,!�`�(i3w¹��<d�Ji�];���w¹��<d�,��L��!�`�(i3n�NQa"_�?���C[u��oŹQ!�`�(i3EfVNN{s�ܱ?'�EfVNN�����1I^�e����kn4@Q�/�!�`�(i3�EhP�Q�ug�%Y��̗0z�cULj� 1��k]m����� ���*�7`����\Z��K���Pxە���!�`�(i3�%=��Lg�%Y��̗0z�cULj� 1��k]m����{"gY*�7`����\Z��K���Pxە����ݚ�Н�[�л���7��{��W�����A@�Q��ǺΕ�A�m�(�]�	��f�?ǉ�=q�\E��0���N��t�3����_�Ξ)�N�ǁ�f�TpD��ZOU	XT�1�wӨj]h�0)xU����V5VM�d|�v�W��I4��欱���j����,X�|H*�ݚ�Н��9+��������i��W��¹���I��RhF�� ��*�C�ժ*)xJe��hy��)]W��7#OOJd֯�y��j��k����U{8�C,0�?���!�`�(i3E�l�����5Ƈ���	I��)���W�w��fD2�e��P���x�NS$x���z*�7`����\Z��K��itXgWZ�G�+5�4��c �&A�5I��RhF��F4#_�h�L�R��k9V��	��y:�^c��D`���J�.�$`b��8�>r&�N������8�C&y8_��s�֙4�(�Ҁч�+5�4��c!�
�!��V5VM�d��0�8k���;_��8W�w��fD���4�-lT��{B�z��z6Y�m@�<����I�?g�f��Qө}�_g�?�H���w�1%`Y��V)�R�7h�,b0V�u�Q�������htO!��nT�Ā���-@��F~*7���&�_���/���l�m��Q�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=Ĉ���rl�خd���!sH�\��X�u��
)\Y����4MT2g�ȨQ�?�Q�_�������� "5�]SƏw0��П�+�
8'���Xw�j�7��9*�"FP��� �mD��.1|��m���tN�w,�������-����rs�i��5O
T������Q��B%��>&ޝ�?1P��+#Cxz!B��[b�0<���:��]]t�GR�D^f�Nd+l�Yҽ֗��J~xAU�"t�{#	�x�z��?�9��V5VM�dn�0�I4��欱���j����u���tt��2��}��M�p}��ϟ��7�4:i�P.j*�7`����\Z��K���t���.`
 ֢����oC���b�J
�g��*�7`����\Z��K���9�u���=3Lv	̅��Tl�������l6�bs��2[������	�;�;b�-�2�3?���*����+7:��a�si՝ӥK�'��iG��Ӆ�+��T����oGo�Z�K����ހ d����M"`h��@�ϸ��#|S������3[�u8�������ET�,/r�UY����7���{r��I`1R�Jʬu�H,qy�W���`moF˯�+)Ƌ��_��F˯�+)��&�C�/n�NQa"_�?���C[u��oŹQ�>b�eIG�5�}�]���p.0��I�!z���.M0��s���4@Q�/�Zt%��m&<	.������Z鎬�������(���ڔ6�.���Vd�2 ٭H�So�x��r��|�\m��sG���MY�{'%s���F����:�#�.��N�x%�M�RG�_`�[4���$[�л���7��{��W�����A@�Q��ǺΕ�A�m�(D}����4��2��}��6d��H�_�ϟ��7�4y��4��U�*�7`����\Z��K�����{�\Z�{k�h�+m��b�;1�#�r��8��vJ�F}��I��RhF��L>�/�G�P�v	��Y4]:C�2Y(���˜V�Q��ǺΕ�A�m�(D}����4۝�hy��)]W��7#OOJd֯̇i�d�?��˺�Q���f�?ǉ�=E�l�����&��Z���,2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!/��KJy����YVctW��X=t��w���'�G��49�V!��#%�/��Z>LW� ���bs_W7�]��m%�/��Z>L%C݇-�%;��|B/B�Â���&S�rD�1�:�Ω�յ�'�)���Ҷt���,iڦKt�iZ]XF�hx��G��!�`�(i3n!��i+�ť�n8���L��g�I��RhF��8usl�z ��ݚ�Н�w¹��<d�Ji�];���w¹��<d�,��L���?�Ho2��O%��<��=�>�t����oD�c=p�J��w x�·���~X�~���$^!�X;p`�����?�dv��oTN֢&@��&��|��p8=�[Ǵ��p���@Z�_F�k-�H��bf�?ǉ�=�|�)՜�4z�Gb��P�!�`�(i3|w�{P^K���3�<�p�� �&���ç�A!�`�(i3�\�!wn�ř�3�<�p�� �&�J�I�'!�`�(i3+�uB;y�3�<F��׿]!�N��y|N�F?P�.!w�E�U�P�)>�
��`�;��%YM�	�v�3�N�ǁ�f�TIX�����^�̷ؠJ��:����_$U���b.����{�vWދ�qc:`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��a���k�_g��������B���+�ϸ�i]T�o8�'��$zө���)󷥯��v
*J�X�$���jh��f�+�t�3���D��m���*�7`����\Z��K���&����$�HN��R��?�d���&��_$U���0�(j��0o�{E}́�9��,'6�F��K�J���1&NXs���ls�uH��q�/���˚����Z��L�{	����F��׿]�v����D�ه4�tZz_nÑ2hꬺ��1�$r�t�}iV��	��y�� �P�qN,t8��og���;_��8W�w��fDbYގEV�9^�o�a�!�`�(i3��;_��8W�w��fD�M߯�Px��|�������x���	R�N~)�j��N�����?�d���&��8�E�"0���a?�5��	}�@�r�<Uee�N�����$��̼�K���Z��L�{	����F��׿]�  ����'Z鎬�������(���[���-��G���۵z �+5�4��c5 H��d��$Ι��o���ls�u!27Ք.+��o������	fd�c�=���L�:w��G$��a��V�K=�u��HN��R��?�d���&��@��i�fKw�R���y��0�J���y�(�\tu2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڧQ����7��� -Q�7�p�D]Ї'G�+R���o��_�Rv�䩲$��8��I�:Fa�7���z��O��Y#&����"sS<�0�zG�������&G;�x'_|~�뽢�7;��1��J�b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-����Dw\����>�lj�Ǎ0Y�{'%s��v�9˞�g��+˘\59:��lJ���l�}0���	��+@f�Nd+l�Yҽ֗��
i#�"��$Ι��o���ls�uGR�	A�"HN��R��bP�63Z�t�5ߧE4��Fr��j������"��Q�JL����	ǜ�N>$m<m��ʘ['Ӭ��yb5]��o�������Z��@?d�s�8K,Q�\C�8�Hj\���n��\��d�٣��c�A�L'�c�Z;�b�R�wX��d=��¾ȼ���4ܱ�������{(z�Sb�f՛ةmy�m���~��Z���Rk��4�����b	��}���Z���7߷M�,���9�ԖY]�蒾�$O�L~�4��>m~�jxBQ%d"Y�9��$9��ճB*�2����CbZ�� Le=mlf�u�c�n��X�L�5_$�՗�(�[�#}�P)-]��h4W�7���\��	���.��yV�$�DK{Eȷ	{�z�� `�*�bn���==g�׷kM�#�> _;��i�1�CɀU��ڞ���ˇ���/�����P��?�N�ޖзu��v�<fGeY�:[d�d���̖b�K/P=<>|�`��c5�J��0�~�G��-�HG($R�i�Yl-����<&Ѳh��N�M��n��mC���!��1{�F}���V6��}�.�p�'�B��?+���נ2�9��V�9!�`�(i3!�`�(i3!�`�(i3̓@?5����T���b�Bϱ�� Q`)��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3/��kOT�)�����m�q�/�Wv�A���U��)���Y;e�iK!���d.O.C�U��B��-����A�;�>��z����8�Hj\�����1:��xjzӝ���I(͂��-����Dw\�����b�S]���o"83�� P�jc�8�Hj\���M7#� �6���n6��dh_��tCdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3G��-�HG($R�i�Yl-ۼ��%�ۙ�b�S]���o"83�C�
���W����Uh1݇S��;�q�Y{�<���^�[�-l��NMm�P˙��b��Bg�Pڹ�ԑ�b�������`y����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끓��~�L ��j�Y{�<����
�9�v�T�T�y�8�Hj\����Fl��m�q�/���e���W�ɸ}(��:)�
�9LeQp�K���&�K�VF�P����9��g�ܧ*ys@B�u�.��.f���s��1�y�n�F�:)�
�9o¶D�ν��jd�	�!�`�(i3!�`�(i3!�`�(i3��j�4�q��_N��¼��=B��u��;���� ���J���*j�B3L���(�Q8;��|B���r�����EHd
0Ki�|2;$�J��7�OT�,��7=���bڕI��.Eqb	��G��W+��W��P����9��g�ܧ*y&tS�D������_�t���׻�fĉ>99��;��|B���J������
H=V��	��y��%����,$�R��aT��3G?�d���&��ҕn�s�[dv�*s?���[`Cw�H���-k��O�)"���.>mT�Ɍ-';��|B�S��sF����b�S]q�6��^�!�`�(i3!�`�(i3��$�\%eK��J�x"V}�IUr��� �&A�5e�J�Pn\�pD��ZOU�S��;�q뽢�7;6ik!�S���{ �4"-�"#+p:wH��|2;$�JأͽgF"?��7=���bڕI��.Eqb	��G��W+��W��>�:| ��k�4eYy�tDWfD.v��W5�!�w(�y?w�R���y�-.�zP&K��Q�m��)� �.�g3Z��~H?��2�.�|�e$S�Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h^·ʌ�C��]���Ҙ�9 �/����P�����
T+Fb%��C��:O�����=�w�����5�O�%E#Py�y�Ż�"�_�0��(����5�?�J�Ń��ɖ�2i�螘c&��,iڦKt�iZ]XF�hx��G��!�`�(i3��иܖ�:�>Xn6��M���o�G�m�?�C��MZt%��m&<9U:����_-�ȩ:[�x�X���+���LQ�f�?ǉ�=Z���ֳ�3�,}�����R8��9$�M�I�h�z�qw ʲ�ݚ�Н�w¹��<d�'��5��s,ݕ����׋�es��O!�`�(i3Ĉ���rl�����@�u��oŹQ2Y��kک����Q��K5���Adu�Bg&��C��[�Do�9�ݚ�Н�8j��zJ�U<�i��W{���铸tC�8�J�Q����q����k��,�:�N�*�x١w��zj�R̶����N�i����b�'Be����s:��i��NU�q�\E��0	ozqP.!ū�ez�,�۞��	�|$�kJ��_F�k-�H��bf�?ǉ�=̇i�d�?��˺�Q���f�?ǉ�=�|�)՜�4�vIn����F?P�.!w'L& �N�	��i�(\{ف(�7���<��Y���U��+�Xa�H(�˕��:�EB�Z5�O�%E#PQS��:Z�7G��#{Ձ�=�niF=�xo�n���㬺����D�Ϩg��U-�e a⣃_B7�}�!��N��	�Ȓ�@{2귑�'=��!���wTR}�/�����y���|����'��$zөI��)���W�w��fD�g�9��,Y:�{]%sշ���⪞mf��EYzȧ���2��'B>&�&i�+#c����nS�3�ǻ��d���!iЈH�����2��C�y��1Q(N��vj��$_.��45��U2X��������,�ǰ��������2܌�I(�g�y��6j�"Hs�l��J�&'L& �N��ƟA#F�Z��E��3?�d���&�P��T�xN���G߽�nh�z:�q�2�_:��p\I��� ��*ȑs;��|Bc^���H�6:�f�]�SK���Bl���O�V��	��y�J8�ȳ4��J\.=e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcKptz�~_%�>�c�
g�[^^�M6Li��.��1�:�Ω�=A���>�LZ*IV���^������)�e��|��x�l��1:�N�*�x^�R@Κ�2���ei�&8�,�뼥<7.���nH�W�f�?ǉ�=Pt�d��R	}�������O9��Q��Q��O�بeD�I��k�+9=�m�n���֣��n��-����� �"��V�E�-�9k|p��z~�I7��-5�B�wj$g�u~xgA�������S3CO��REԔ	�8�����ϲ������i���i�\�>&�&i��&�C�/W����vcy��<
DN��X;p`��d�uY�ؤ��E�����|>U����z~�B�wj$g|�����ݪ���k�+9=�A�����y������i�-�����m l�o֭�B������t��˳3[�u8����ꀍ�U젩`#�4>?� �1Y��
�iC-����b=���
�	?�<�&8�,�g�Hn7�(�?V��j�c>ݣK�6<oC7z��R���V��"���q�rVu,� ��u��g��L�����.!ū�ez�,�۞��	�rVu,� �+��%�k<�6��w�6Y����$��%�]�
�R��];�1�+ptA-I�p��g���^u�� 
~�F�,���XF:������X`��w{���Z���F%�X��O�_�-��0��ԡ�/$a��F˯�+)Ƒॉ,����g��U-�e a⣃_B7�}�!���:�,���P�,'",H� ��ˀч~&5�r|�g�ܧ*y�Y#	߾u}�	76�&�;��|B`#���J��M�r�!��X�.����2܌�h,\�NyVX��-|?��Vx�%Ls�N
�u�}�T�\ ��;��|Bc^���HV;ƘdO��cb>�h�D���b8IU_h�¦�naä��,bxqX�����,�ǰ��������2܌�I(�g�y��6j�"Hs�l��J�&b���J�/�#2fک��HC�d��g�逑�D���H��<�C�Ar��� ����Dɵ�p�AJ�e�$�X`��w{���Z���F%�X��p����*EYzȧ^0ػ]Yt�Y�7#�xI�d5z�R��T�\ ��;��|B���r������f
t斃�B�ӗ�zjJrf����G�m���*J�X�$����q(	�fw�R���ykb>���p�JM����&UX�{6j�"Hs�l��J�&b���J�/����+��te��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc
M����n���2�V��cb�P����T�}ɻ���}J�|���|���/Q�������d���!iT���/A��'HY-��Yk"1/]���!E���VG%�z�y�l�&�����S���� "5�]9��n�7�Y�9ηd��K(��-�f뼥<7.��H�ʱˡFZd6�o��zg��p��I7��-5]�j}�_U��TP���D1�Z���=�,���9^-�x�	�2��GF��a�1�Z���=��o�� ������it	�TU����z~���MK�LS�_�p���it	�T�=��?����d]���g�P�e�9�y�3�A�e����kn4@Q�/�!�`�(i3���ꀍ�U젩`#�4>?� �13Lv	̅��!�`�(i3���*[UxG!�`�(i3�չ�Ad���c�����:��IK��<EOJ�uxm�3���w�@V�?ZFw�Ns+��6�.7��m�K�!�`�(i3\.�l���/*;63��dn��A�v���{	���Dv��Y2\V��rU�w�⽒��8�>r&��H�ʱˡj�:�IL;��|B�6�����O�X�aY���	��#<�Eg��ߘ�)�I����D�Ϩg��U-�e a⣃_B ;�|4 w�A��AC�m;��krk��+�� mч~&5�r|��u�)���'��$zө�Ձ�B#�~;��|Bɖ!v��Z�
�且�.�g3ZE��g�Hb�t]�<Lz��al���Z��E��3?�d���&��q@�?��� �l���hu*_��� ���J2��������������T���Ӫ!�J��:������*�t��v+�/;$�������1�1F%јI��/z*x�n;��|B���O8k�Ĥ;-](�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�u��Hic�{0��d#\� �6���B�@o��[ea�8����U��}�o���#��X�����S���� "5�]W���`moF˯�+)��h�\ƙk����p�><��d5�:�w�+���LQ�f�?ǉ�=h�5,Wlr�r%)cANU�:|��?�R��n���Lr�VU����*
��c�<v���G?d��A ��+���LQ�f�?ǉ�=��h;e��w���U���І��%n3uZ�v|�E��n^���+qѭ�+g[���|��pe���b��˺�Q���f�?ǉ�=k/�z�xEQ�苇��Fe#OOJd֯�|�)՜�4-��r��gGr�����rk���6���
|j	FQ�)HVi�p"���#?�q�\E��0M7$����1Ʌ�Mi��������<�ry^�$���]׽��X;p`��D�����M�;��i_2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��"/���]�Q诤�e��C�`�/�t��cm�@�ᩖ%�!����5��fH�6J)�s���-�)��|���=f�}��U�����̾0���;���˔����vg�ĝ����a��X`��_/��;�y/Ә���@�ۻ|2���̂; ,@�� د<�l雲�fb�����m� D�@G��l��3\s��$�Z;��|Bc^���HP�a��t�'����9|s��^<4mB�@o��[�|�hJe�A>��*�X�3�z?Z��ϸ��#|S������3[�u8��� ��w��]n���І��%n3������k�+9=���(��U��֜��3�AQ�0G�C�`�/�t��ߖ Y��U���gFck
�������}g�2Y��kک����n|�p[Y���"����)�-}�|ݔ�3�z���.Mp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���K+!q���!�`�(i3扈�[-�c]^�mOeTky��2��}���zgm##�+��%�k<�^�V��	��y�3�&A��SwE�=p��-:�N�Ò�}kutC������i{��*ȑs;��|B�Տ� �*��q�)�`C�G����]'\gWg��	�Z�kfc?�#	*]]�(&�L�xjzӝ���I(͂��-�����2��}��cVe�U2�<��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�G`B� �'����u��r���2��}��cVe�U2�< 'J��@�D`ks�F⽉��%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}���Q���!���ūaT��3G?�d���&�s͟;)f���KXL6�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9Y���&���'܍|Cy���QJ�wk����\����|ݔ�3�(n�'�(�S��)��R�^Ƒ��;��|BEΟ��
�U�a�(��^GѬ�_���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3�v�Wס���G�K$x/��&���PC-��i0Q�͹�Ɩ,�b�R؅�!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3��Ě�����}Dq�f��3��C���H�� �YߥթD�[*�Bi�v�V���;AD�e�{�W!�`�(i32+5�"�����-P��F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊<���He�ylB��-t���m�� �ݪ�򈟕��+�v�7��]�ݚ�Н�3��0����g����F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊����xQ�e�ylB��-t���m�� �ݪ�򈟕��+�v��t���?�� h�ҩ�!�`�(i3�lTN��I���q�}���{BO���5�%]���a(􆿳����^��!�`�(i3��jVѭ@!�`�(i3u?�:�H�jsrCm�k�J��6�d�t��w��X�'����u��r��!�`�(i3q�\E��0��@Z���rs�i�}�O��LTSG��ʎ�=U9��R�^Ƒ�Ӆ��I�ѪtR�^Ƒ�ӆ�v�9��!�`�(i3�����!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1��#ƌ/B�ݪ��2�r5�����jV�{+�fbmDF�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ o�n�J-�ƪe�0c�)�Ul����,�ǰ	r�R��Z����i�|7��_	�s�t�{���6������]'m���G�K$xE�p4rqG7]u��
�3�R�^Ƒ��;��|BEΟ��
�U�a�(��$��,Ix�6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^q�\E��0��@Z���rs�i�@24b��H�[���wkL�1p/-��G�<6�U����z~)���	6�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=��X�z��V��	��y�߬9�6ש�ڔ*��T�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc
M����n��i���~+�lX҉ޖ�˞,cƶ��^�}���8�\�(fw���I��RhF��0��N�F�6��9I�u��'����(fw���I��RhF���,�=R�/��Se����-���^��U���P[�񁫴}2��uR�9$��i����t�T��?E-h��`f���sC>��Ӛ��S�J\7!c�2���j"�²O�y���0ܔ��'ž1�|�'����u��r��N��r8!�k]m��Z�����hh��,��Oˊ��C����t�ǊS�>�!/�_�n�To�[
MQ9�F�1�m+�D8�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*�Va�ir���M��2"���&�^��v�8:?�'��ᦾ�;���8���U�._�nQ�rV��q�t7�v�]��1���U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^N��r8!�k]m��Z�����h���G��S:t�L)��k]m���E��Y�^�Mi~_�T���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�������c����g��U�S��q�}��il���iA'R�	z�#,gB��Pߺ0��A���ۖ�)�-�W���a�x�G9�:Q��Ĵ��ޯi���l`Zd�g()��ikp���H�����[��l_G9�:Q����v�z`���ө%�Sg()��ikp���H���׾ŞWsuz��"]c�#y�>�)L����0ˮR�m ޶&�hbvk~�#x��#�H��+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!H�x�7X�J�����_�U*Cw�Hm���9��N	{8G9�:Q��Ĵ��ޯi�I#�(���)x�?{���x.�Knq^nї�Y�_�n�To�[
MQ9�F�����
��\�H��/Sg�w��'o�v��؄aX��I�_Pg<�l��姹���Mt��a�x�]c
j���l��姹�ȃT����A���ۖ��S�<Ԣ������f�l��=5;֡Q��Ⱥ���>��� ӫ/��m�D�K��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6��J�����_�U*Cw�Hm��G9�:Q��Ĵ��ޯiڼ�ze��>տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<�%��g:�����<�ׅ��A5W��v�8:Tr�E	�[��J�����_�U*��ө%�Sg()��ikp���H���^?������X��O���r����!�`�(i3!�`�(i3!�`�(i3�I�_Pg<�%��g:�����<�ׅ��A5W��v�8:C��4�I[��I))����A�m�(�-4�{>��G9�:Q����v�z`�Cw�Hm��G9�:Q����v�z`���ө%�Sg()��ikp���H���GM��QО#y�>�)L�/|w~S."��*Ha���J*�Rs�0��|�_�Y�j�W��� D�cg�}��m���+)x�?{���<m�N=-�w���+ާ�����ݚ�Н�!�`�(i3!�`�(i3 #��zG���J����k̇���APߺ0��A���ۖ�èr�L��b��v݋N�����&r�"A��A���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~��0Ր�5Ҹ�u�����φ��<�6�@a� ��fFMqlgd�G}%����3fUi���Z�͗�M9f��;�jmT�#bs��2[�a��o���H�RtV�^�}��il��o\�B/�k9a�S6��_
�u �V.��$��l��=5;r�$�(��{�R���/�O��� ӫ/��m8D����#U��,H/���k��^�1��dc�@c�����h��-����;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�j4�����ݚ�Н�޼QE1��v1a{J�)�H�b�b�Bϱ�G9�:Q����v�z`���+_AdV
�:qEp�;�P�t�5fĉ>99��A0ok�׹��*P�{���"��\��}g��V�;ܬo>v<~<�=a��0� ޼QE1������m�(��k8!�`�(i3!�`�(i3!�`�(i3!�`�(i3+�F�$-�S:t�L)��k]m��l��e b6vJ�pZ� 4�F�Α��Dr�2�N��r8!�E��Y��Q�
w�8D�t�%o�V���-$�!�`�(i3!�`�(i3q����`U�0�V;�M�J�����_�U*���$����;-�]�pR�$5iL�Pf8e���N��r8!�E��Y��Q�
w�8D�t�%o�V�g�yl��6T�T�D��ao.\C�k����S�{؁C�*&#�4?�o�5�h�B�c\��L̎C��fx'v�ao.\C�k*h�!<^Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������Mڷ���o\�B/�i
�i�w�Qטg�u2�Tt$Ó6N��o\�B/7� :(c�Wh<�!C���>��� ӫ/��mo��7�^�1n��y��a3G7```+��)_�32�K�y؄@�!�`�(i3!�`�(i3����&��+�%�t�*#y�>�)L��H"҆>X������*fW� �/88n
I��jÇ+�_�n�To�[
MQ9�F��,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcU�۩}�w��k]m��
ae���K�9�*��� c(H޵D7W�:���iޚuq6p��j����Q�9�|`ЉɁmwlc(H޵D7W�:���k!��,�<��y�@�v,����.�u-�w���+kGA��ݼ��r����!�`�(i3�o�5��!<��y�@�vFn�H�~M������f�l��=5;O�R'o��!�`�(i3sU�@{Q�p��j����Q�9�|`ЉɁmwlc(H޵D7W�:���k!��,�<��y�@�v,����.�u-�w���+�\#���Ƹ���r����!�`�(i3���>�t�mo5i,�Ĕi��)��ۺ��fyd�,m �\��\�H��/Sg�w��'o�'uFէ���p��j�����8"c�։Ɂmwl�E��Y��Q�
w�8D�t�%o�V\�Z�0��9$��i�Yi䚠疛!wFii���_�?2��HL�U���W�H�2^�/3!�`�(i3�0�9&،�d�G`5[��{#Ÿ�&Sq�a"��ř�!�`�(i3!�`�(i3!�`�(i3�����wP?��i/R�c��;=~. .����mo5i,�Ĕi��)��ۺ��fyd뉯ӌ$/k�&U;��]�x�'��x!5�kz���[h�x�1W0�-��4��Ɂmwl�E��Y��Q�
w�8D�t�%o�V�g�yl��6T�T�D��ao.\C�kT���/T$�&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N�����U-�pë��";Yy\'{w#/ B!�`�(i3޼QE1�&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N������G������p8�Iט��ō�Zm\�l��ì�A؁C�*&#�4?�o�5�h�B�]�{����d�G`5[��{#Ÿ�&Sq�aM^�ؾiZ-�w���+�gVdxQ,��a�vw����~m�(��k8w��?L�@���wp>�\�H��/Sg��'|F��d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[���&YH��-��k���H�2^�/3!�`�(i33��0��e��0�U+�qbp@��C�7ª6�9$��i�Yi䚠�5���u�L�!�`�(i3!�`�(i3!�`�(i3��c���鿉�X+�kQ��v1a{J�i�\��ou#���3qV�[�U�b(l�rD��ЀUg]�6��;b؁C�*&#�4?�o�5�h�B� ި�6v ӫ/��m�h��"��^����'5��9$��i�Yi䚠�@CF���(�b��v݋N�����&r�"A��ArS����u�}�Q���GM�о٫�S��wE\�!�`�(i3!�`�(i3�I����~u͘6��q���j�W���]�B� ��8@��1�*)�2�"��wb���E�¸>`!�9wY����<��y�@�v�&Sq�aj(��;����_��%$>_�n�To�[�pI�
KrS����u�}�Q���GM�о٫���^O�K����fx'v�ao.\C�k*h�!<^Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������Mڷ��iA'R�	��}E-��$@PJ+5*�轓�A1�J�����_�U*����e��ھC��'#���fx'v�ao.\C�k C�Mh�n �O`�Ag��ۭXX�|ʡi�����Fz�!�`�(i3!�`�(i3����&��+�%�t�*#y�>�)L��Bѭ�pR�$5iL�$�F�V��&|���BY��l��=5; �e� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���Mڷ��iA'R�	��}E-��${`�9$��i�Yi䚠��&���)"r�DyA�S⏸[����LG��&��a�vw����~m�(��k8���wp>�\�H��/Sg��'|F��d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[���&YH�HL�U���W�H�2^�/3!�`�(i3�0�9&،�d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[��H	X�ʁ���Mյ��#�@����ۭXX���E��O��d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[B���v��؁C�*&#�4?�o�5�h�B� ި�6v ӫ/��m����	���γ~<�����6Bj�!�`�(i39<��`f;]MBg2Zr�G� Y� {l��	z�9^Ȑ�I))����A�m�(�W[����p8�Iט��ō�Zm\�l��ì�A���V��H?Ә�%"Q�ܦfM� �'9�5���c(H޵D7W�:����p�A�ԍ'8�����";Yy\'{w#/ B!�`�(i3޼QE1������m�(��k8һ��6�!�`�(i3!�`�(i3!�`�(i3�����9�Xy+�Mk��趵��1�F���������m�(��k8һ��6�D��)��	u�}�Q���GM�о٫��s�~�L�1{&��� )S���z;]MBg2Zr�G� Y� {l��	�g�yl��6T�T�D��ao.\C�kT���/T$ǩ����m�(��k8һ��6ݕ��wp>�\�H��/Sg�u-Y2�G�1{&��� ���xl�ݚ�Н�!�`�(i3�V3���L�瞩w�j���@ΙN�[���-ل9�#c�ᜂl��=5;J5�#Z�"r�DyA�S⏸[��t��7�M~�V3���L�瞩w�j���@ΙN���HPԎ��V��H?Ә�%"Q�ܦfM� ��x�1W0�-��4��Ɂmwlc(H޵D7W�:����p�A�z;#o"�I0���ԏ�ʖ�:���V3���L�瞩w�j���@ΙN�[���-ل9�#c�ᜂl��=5;� Ek�0��������mo��jVѭ@!�`�(i3��dN���ub�z'hۉ)��_�2��|2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��7&���Y'=�t%�!�XH��Oi�HU5��)4�3Yb�J+c%F���_�z<���L1v�}7>�W��	2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��:�dy�v1a{J����%]+a���G����E������7D!��l��姹�xAQ�Y;x����̜�I0���ԏ�.fOe	���X�a1p��j����Q�9�|`Ю�K49AԢ�a\�[�U�b(lƿWdM4@��z(��xo}E�٦���sC宸I))����A�m�(�QNȮ���k/��m#ׇӭ��!�`�(i3!�`�(i3h큈��{��UJ����"]c�#y�>�)L��H"҆>X�(JdT�ݙڈ�KK?B�&�_j����)Ł�I��jÇ+�_�n�To�[
MQ9�F��(��&��[��m�U����#34�?��˧+P"G�wk�[�S��]c
j���l��姹�I�oൠ��ڈ�KK?B�&�_j�In)0LH�* �b�p�Ĵ��ޯi�-Qq��Pn���G��(��{�O�iA'R�	��}E-�c��n�#&|���BY��l��=5;\�Z���O`�Ag��ۭXX�|ʡi������ڈ�KK?Ba���$_Ĵ��ޯiڡ�F1�4WM7�FM\�1�����\�H��/Sg�w��'oª���#oMA�H4$B����>��� ӫ/��mt�����W�br�*7�iA'R�	��}E-��0��ٟ�͘6��q���j�W����+G��ܻ�ߣA����Dr�2��c���ğ�%��g:���
A�%�q����	�����͘6��q���j�W���]�B� ��8@��1�*)�2�"��wb����,]�������ڈ�KK?BD�1N��λ�g��ZR�,��9 �ubK���E�g��ZR����z�Ji��1ʟÛm�w��ГQ�H���&�b �hvT�+]�x}NI0���ԏ�.fOe	-=3�$��ϐa�x�����on�b�Bϱ�m�(��k8����~�䱢�z
A��Φ�gz(AٸI))����A�m�(JX��!�.�`;���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq�(Ul��?U�D�K�X�K{�(��	}�@�r�<Uee�N�����b��[cS;��|B�V���p�e�S��@��Vd�uҹW3�"b!�`�(i3!�`�(i3�s���6�v1a{J�o1J����٣�}��iA'R�	�z�?��D@N�ǁ�f�TpD��ZOU���Gx5��WdM4@��_�U*�>=:9_�aV��	��y���x.0��X��FO��(���*�`�
��pF泥���k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��L}c��ko#k��^)�Qטg�u2�Tt$Ó6N��o\�B/�&���+��h<�!C���>��� ӫ/��m�D�K��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6�JeYSWe^E1��b���S�C���0�V;�M�J����'",��X��a�x��"�%�U_k���$,@����:_��k]m��Cw�Hm���V3����C��z��&���)"r�DyA�c(H޵D�ҏ@n�k!��,�Sc��h� ����r-�w���+kGA��ݼ��r����!�`�(i3!�`�(i3�V3����C��z�ob.�Y�2W�b��v݋N�����&r�"A��A���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~�z5�0P�ġ��x���u�Y�KG�ξ���I��RhF��F4#_�h���Se���7�}�!���e�S��@��Vd�Y���DO�!�`�(i3!�`�(i3a�u��e�MN*�������*y}e���:�#�|$.@L�`f�Nd+l�Yҽ֗�51����~�gKh���V�H�M�I��)���W�w��fDl2����}*�NRcnvyw�R���yW�R�w���L�>5�C��Ҁ"���`Vk�d��f�Nd+l�Yҽ֗�X�e��n�ސ����U��)���Y;e�iK!���d.���+�^n=\f�5>�HҰ±�͹�uR�:l��xjzӝ���I(͂��-����.[�Kδ9����˦G�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н��I��� g~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�P�궊�2�����8!��?V�ы�(�)x�?{���x.�Knq'ێ����� h�ҩ���6��5=��)Q��h�xF墣c#���K!�`�(i3�����!�`�(i3Zi=���lr�{��|e��0�U+�qbp@�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�d�n�ͻ���~͏닓.�`�3���M��,�IX0F�MV�ҁGG%4vkz����`���φ��<�6�닓.�`�3�P���F\xjzӝ���I(͂��-��������FYs%?es� e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3<�g��H��&�2���)x�?{���x.�Knq��5+*��d�@���G�X���.��ġ��,��5+*��4br���qP�V>t'�̗����S]�_�_��u��r��`
 ֢���֦�n��{_8�Y��=�}�Vݨ��}Dq�f������!�`�(i3s�3r<��AgC�&��������5�,D|r9�g()��ikp���H����m-F���T�YN
��)e���T���b�Bϱ�h�5,Wlr�r%)cA�5QN���d>�c�n�P3�K��b� h�ҩ���6��ZRR����Mn__���q�Ӯ�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MI8�ѐv2Q{VcҟA��0Ր�5��v/�(%줄$�HY�����A$�P������5d��n4s1�U��B��-�*P�{��Ɖ�<�(]|kY-�xjzӝ���I(͂��-����N��r8!S⏸[�nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��u?�:�H���^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���Fie6ӭkk�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н�޼QE1����"���dN�<@Iv��nt=:��:5A��p��w�w:�!�`�(i3^()��>�����U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^M�yx�,�G��i/R�c�${`G7```+��T�TN��!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M��uR3��%<�X1H�w���ސ����U��)���Y;e�iK!���d.���+�^n=\f�5>���u����uR�:l��xjzӝ���I(͂��-������T��xW����˦G����P�|T�T�����U(���B����Ӝ$��BS�>�!/�_�n�To�[
MQ9�F���v�9������g�Z��3��a���!@�f")u��r��܌;���'����u��r��u?�:�H���^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���Fie6ӭkk�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н����cJ�C����o�W�F}���V6w��EO"�̞��>�_9�R�5;�/�O��� ӫ/��m�QP�*Hd��:5A��p��w�w:�!�`�(i3"G���RG7```+�ֶ������YN
��)e�W�J��H����8�O�5���1tSjv�!�`�(i3pR�$5iL̻��Fd]�ob.�Y�2W��C�Y�\�fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹��Li�AE��� �Rɴ��S��)�5���sO�v(�y��U��)���Y;e�iK!���d.���+�^n=\f�5>��UE�'���(0̈��N����"sS<�0�zG�������&G #��zG���J�����/t4�q���o�F}���V6� ��=y�̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q����Z$�x$�֯� W(���27:։�X+�kQ��v1a{J����nFy� �ֿ�JO���%>�rGO�D mWN��Ě���aT��3G�IX0F�MG9�:Q����D����1����ciAG9�:Q���O7�4[i�$R�nS�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2���j"�²O�i.����bs��2[�a��o���H�RtV�^G9�:Q��Y����(��U� �,\���͔5��:m�\�H��/Sg޶��"���̺`����1�����\�H��/Sg޶��j�}a�cfn��ٙ��Z*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81-���7,D|r9�g()��ikp���H����m-F���T�T�n��a��#�GWW�<om���m-F���T�YN
��)e�W�J��H����8�O�5���1tSjv� #��zG���J����0;�������G1=��͘6��q���j�W����΂o����^�?��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxģ��_�ڑ8�`Lv�RU��P��i�u�}��il��J��O�����!�o��_�Rv�䩲$��8��I�:Fa�7���W"�P�K�0_f��3%�~eG���A(�c���_G��Hb� h�ҩ��I�_Pg<�(y�.
جHR��o�W�,\���͔5��:m�\�H��/Sg޶���W�Z[��MQ�'���1�����\�H��/Sg޶��j�}a�cfn��ٙ��Z*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81-���7,D|r9�g()��ikp���H����m-F���T�T�n��a��#�GWW�<om���m-F���T�YN
��)e�W�J��H����8�O�5���1tSjv� #��zG���J�������ߧj@Q�����&��"]c�#y�>�)L�^b٫
z�(;-ob���;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��I�_Pg<��4���Lo�h:E�,�do2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q����Z$�x�vG��*Ha���J*�Rs�0�ǳ7��y.��c���鿉�X+�kQ��v1a{J����nFy� =�r��J*�Rs�08�b(��g]�6��;b#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#xo�������Qטg�u2]c
j�����7�*w#;���W��m ޶&�hbvk~�#x��#�H�޼QE1��v1a{J�Bz��s�V��m���+)x�?{��
0#`�1��׾ŞWsuz��"]c�#y�>�)L�^b٫
z�s�ť���)x�?{���x.�Knqo���n[�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��I�_Pg<�4���TS3���/k��1x�a��2e�>���x��j�W�����ד*(�os}�&à��b��v݋N������M}Ĭ���.�f���I�J*�Rs�08�b(�����̜�I0���ԏ�.fOe	m���h��v��؄aX��I�_Pg<���7�*w��D��q��S�C���+�%�t�*#y�>�)L�b�@_	��)�p��ZI0���ԏ�.fOe	m���h���s��訌��v�8:������fI��jÇ+�_�n�To�[r��}k:�%��H�7���|ss�j�W���yͧT���E"����5�W9a�Fc��Ǔ��K��v1a{J��¸�k�L�����f�l��=5;R�ˊ	18��X��g()��ikp���H�����V1G�׊�b��v݋N������M}Ĭ���E�����{��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6��J�����/t4"����5�W�����G�v1a{J����nFy� �_Y��t��3
�v�v-}�	mpÊ�����j�W�����ד*(�E��W�u&�Pߺ0��A���ۖ禡�Q���#y�>�)L�����/s=s��4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J�����/t4��UH���4տ�:
hbvk~�#x����I0���ԏ�.fOe	m���h��g]�6��;b#y�>�)L�b�@_	�"����5�W�����G�v1a{J���Ꭓ�[���ө%�Sg()��ikp���H���GM��QО#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#xa��H9��k]m����\�6��_Y��t��3
�v�v-}�	mp�dA�M}.F!��D�����k$ !�`�(i3!�`�(i3!�`�(i3�}��il��A�{�>�� ��
�m���+)x�?{��
0#`�1�������f�l��=5;R�ˊ	18��[	�"~�}��il��Rm�㭼�S}�S��� �~�^#y�>�)L�^b٫
zܫ5u�q��	�����aq��uG�բnG9�:Q��F��P�?��4�+��_��A5W��v�8:Tr�E	�[��J�������ߧj@Q�_Y��t��3
�v�v-}�	mp�dA�M}.F!��D�����k$ !�`�(i3!�`�(i3!�`�(i3�}��il��Rm�㭼�A�!�[��5�*Ha���J*�Rs�0K=X���d���fx'v�ao.\C�k�ף�D�~����Jϑ��+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�؈G�j��m&����T��Ŗծ��7W�:��e���b�!�`�(i3!�`�(i3!�`�(i3q����`U�0�V;�M�J����0;����0
"8�'o�*)�2�"��wb���E�¸>`!�}��il��G����1�E�AvY�5�h�B��A�	���\!�`�(i3!�`�(i3�I����~u͘6��q���j�W�����ד*(��j�Y|��a�x����r͖���"��Id�fPa[��I�_Pg<˃�B�1Yw�Yi䚠疛!wFii�"�/̯��3�{s��ֹ圂�Zd��(̚N�:R�j�W���<�'��V�I�'��x!5�kz���[h�\�n��I0���ԏ�.fOe	m���h���,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��L[��m�U/|w~S."��i�*O����Qטg�u2R� [�'a,�v1a{J���Ꭓ�[��[�V�+�6f6,�#�I))����A�m�(};l�-����!cI͸I))����A�m�(};l�-��?�%�'^ȴp��j����Q�9�|`��Y�m�k?j!�`�(i3!�`�(i3!�`�(i3|0u�ښF���A�k]m��5L5@�m��B��رzh4�+7{�R����� ӫ/��m�A0`��A�"��(ޅ���>��� ӫ/��m�A0`��A���/j)	 ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���Mڷ���o\�B/N�.�L�0Ϩ �~�^m&����T��Ŗծ��7W�:���iޚuq6p��j����Q�9�|`ЉɁmwl�F��M:J�5���d��!�1G9�:Q��HN�YH8x|?Ә�%"Q�t�ч�����mo��jVѭ@!�`�(i3�� 3�m&����T��Ŗծ��7W�:���rL��7�_�n�To�[r��}k:�>�hy�!�`�(i3�ݓ�W���"r�DyA�S⏸[����LG��&G9�:Q��HN�YH8x|?Ә�%"Q��(�K��F��M:J�5��,����.�u-�w���+�\#���Ƹ���r����!�`�(i3�VR��)Đ�G����1�E�AvY�5�h�B�͞_'Bi��fx'v�ao.\C�k�ף�D�~�ڭRyԍ���#�@����ۭXX�WŚl��E�j�W���<�'��V�I�'��x!5�kz���[h'9�5���)�5���sO���%�$�m�(��k8w��?L�@^?���W��j�[O����k$ !�`�(i3�}��il��G����1�E�AvY�5�h�B��A�	���\!�`�(i3(*�O�q�@��i)&
�k�����oT`kz��{V�-_8���G�7W�:��G�z㤧{�>
�eEQZ�G����1�E�AvY�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR��M��e��)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��^?���W��j�[O����k$ !�`�(i3�}��il��G����1�E�AvY�5�h�B�$5z&�D���ME�R�, &ấ<b�(*�O�q�@��i)&
�k�����oT`kz��{V�-_8���G�7W�:��G�z㤧{�>
�eEQZ�G����1�E�AvY�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR��M��e��)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��^?����8������k$ !�`�(i3�~�7p����nt=:�+�_0c �I	�����g[�s6{޴�i��)���1�#��d_!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Y���g��{�6G�a�x����r͖�k���$,�C�7ª6�L_v,<=��}�I����&Sq�aQ�y�QF��fK�Ěk.!�`�(i3^����'5�L_v,<=��}�I���Fn�H�~M�y�)w��W�l��=5;R�ˊ	18��[	�"~�qi4�747B��[�<?Ә�%"Q�ܦfM� �L�Y}śT�!�`�(i3!�`�(i3+�F�$-�S:t�L)��k]m����DބiMb�R�f��a��;���=����qFz�}o*o޼QE1�Bz��s�V�r�G� Y� {l��	�g�yl��6�����������iv�!�jT7|�`\%��u7W�:����p�Ǎ�͚�3�_�n�To�[r��}k:�b�	.�� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ht)PjL��k]m���E��Y�"����5�W9a�Fc���F���A�k]m����\�6����~�	hnp�����b��v݋N������M}Ĭ�����V1G�׊�b��v݋N������M}Ĭ���N��E�Q�>�H�(�#ve
��e����R,�!�`�(i3!�`�(i3!�`�(i3��+�t2�a1�����G9�:Q��F��P�?�?$٭n�rD��ЀU�r`�JtоI0���ԏ�.fOe	m���h�����̜�I0���ԏ�.fOe	m���h��֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@��_�U*�^�?�9�*��� ��\�6��#P��Ѐ�N�w�qX�f��EJ,�G7```+�
�HYF�@�����4R�ت����¿'��x!5�kz���[h����XzRL��MWX��\�6��#P��Ѐ�5�h�B��ME�R�, ��Ѻ��	�1{&��� ���xl�ݚ�Н�!�`�(i3I	�����g[�s6{޴�i��)���!D������eW�d/=me�%b\%sU�@{Q�p��j����Q�9�|`ЉɁmwl��\�6��#P��Ѐ�5�h�B��ME�R�, m��
~�B�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\����oW�l0����'{w#/ B!�`�(i3l�[K��K8��DބiML�瞩w�j���@ΙN�z�}��b��v݋N������M}Ĭ���N��E�p8�Iט��ō�Zm\�l��ì�A�����5qo��o�����&Sq�ae:rmv�H�!�jT7|�`\%��u7W�:����p�A�ԍ'8�����";Yy\'{w#/ B!�`�(i3޼QE1�Bz��s�V�r�G� Y� {l��	���-$�!�`�(i3!�`�(i3�����9�Xy+�Mk��趵��1�F����Bz��s�V�r�G� Y� {l��	\�Z�0��)��%��+b�O~1��GM�о٫��s�~�L�1{&��� )S���z�R(R�X���Ǹ���m�(��k8һ��6��b��QM!Ϊu��U)�Fx�Ǻ^U�:Q��z�˔ �y=k�2�u���e�՝*U��eW�d/=F�[$��<���H1���~!�`�(i3N��r8!��DބiML�瞩w�j���@ΙN�[���-ل�{s��ֹ�Em��r�~�����wP?��i/R�c��;=~.T"O5�`�7B��[�<?Ә�%"Q�ܦfM� �'9�5�����DބiML�瞩w�j���@ΙNVB=�4�S�-��k��[�����������5qo��o�����&Sq�aj(��;���Q�y�QF�靰v j}�!�jT7|�`\%��u7W�:����p�AE2p��Fȯ+3�YE\����oW�l0����'{w#/ B!�`�(i3i��r�+�<�W�.�P�@���?���"'�nH/#���J�ďx'��I�`�
��pFC�R��<:�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcU�H8����2[QvA��֣T�5��$@PJ+5*�轓�A1�J�������ߧj@Q�h�%��?Q_�n�To�[r��}k:1x����̓@?5���嚚3�%�I))����A�m�(};l�-������l�Y;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��0<�$#y�>�)L�^b٫
zܫ5u�q��ҏ@n�$@PJ+5S:t�L)��k]m����DބiM��pqo�}�;-�]�̓@?5��l�ҵ�_�k]m���^�?�9�*��� �k]m����DބiM�YG5`FFB5=��)Q�n��y��a3�J�������ߧj@Q�_Y��t����M���X]c
j���(y�.
جH��O��U
h�07�;|''ZT��*�/4{+�x<�;���jVѭ@!�`�(i3!�`�(i3M�yx�,�G#y�>�)L�^b٫
zܫ5u�q��ҏ@n�rL��7�_�n�To�[r��}k:�b�	.��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �b��D�씴SZ���U��)���Y;e�iK!���d.���+�^n=\f�5>�Ml`�`\Ձ���� \���F�`yx�>�+X�M?��y�Dw\����.m��K�+���w�c�c������_
�u϶=f�'�1�����\�H��/Sg޶��j�}a�cf�Lͷw���]�x}NI0���ԏ�.fOe	m���h���%@{Ex���k��^�1��dc�@c�����h��-�����s�Yls��8��GMm�HxX����U�._�3
�v�v-}�	mp
���U{���8^��hJL��;���N�4��N	�7q������O�޳!?�R��nścp�B��-/a8V�Ո���m�q�/��v1a{J��a`p�W�8��b�Bϱ���j�4��k]m����,^�V�:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxMl`�`\[�H�l�b��D�/�����	^%�R���m���+)x�?{��
0#`�1��9a�Fc�����^dE��C�x!�H��SW]#��5�m ޶&�hbvk~�#x��#�H����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcx�dŕ�n��.m��K�+���w�32��B��Qטg�u2c&��n��C�x!�H����'^_J���"~6���aq������n}L�I))����A�m�(};l�-����!cI͸I))����A�m�(};l�-������l�Y;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���j�4��k]m����,^�VC&��b��Ɔ ���Ve��˅���ө%�Sg()��ikp���H���>��B�K�.m��K�+���w�?�H$~��	�����aq��[��n;�D/�����	^%�R���m���+)x�?{���<m�N=���fT��F*�L��!�`�(i3!�`�(i3!�`�(i3;�x'_|~� �S���}�cЉ�M�+!�j�8�3
�v�v-}�	mpl�!����_�n�To�[r��}k:�b�	.��=��5a�y�iA'R�	:�@�F���,�
�CA_�G��-�HG(�b�'BelĈ�\פ��
y���)_�32����r����!�`�(i3!�`�(i3!�`�(i3�G%�MP3ö�3���:b׻���3�v1a{J��bC�����'�NKc�F�*3��ö�3������7�V�k]m��d�r����dQ"��؆��)x���l��姹�-��#��e�S��@��Vd�2 ٭H�So	.���T`A�WdM4@��_�U*:J����#SX>tG�zi�X�+2�ꎷĬj����M��v�}졞���$U������h�̯#DC���C��Wo9����4~��E���ZaL݊���2�"�G�p�Pڹ��/^�w?�d���&���5�G
m�D ML:�N�2	�����8�5�IX0F�MV�ҁGG`5:�����+�^n=\f�5>����5��M������S������"sS<�0�zG�������&G��6���2[QvA�΁�a�n���I����~uK7͍��|��W&":�ݚ�Н����D)�ܮ�S�Gz�J�a$�Y dN�<@Iv��nt=:��:5A��p[�t��#��l��姹�g�YӅ:�E�g�������(ӈ���m�r����١w��zj�v1a{J�&��	�>�n��>�my$�N��o�/���;�/��@���WdM4@�k̇���A�C��|uK7͍��|��W&":�ݚ�Н�K�\7}�W,��+G�����̑:�dN�<@Iv��nt=:��:5A��p�T�T�y�/������Z� ��(HE�g�������(ӈ���m�r����ЈH�����b�'Be΁�a�n��n��>�my$�N��o�/���;��6�����
y��!�`�(i3�I����~uK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv���6���2[QvA�΁�a�n���I����~uAԢ�a\蟴���P`��ɠD(c!)��w�K��r�]�4�P�l��=5;���o�1g��U-�e1�S�������6���2[QvA�LO�>��
�I����~uAԢ�a\蟴���P`��ʱ�O��W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3�⒍~����v�z`�!�`�(i3���G��(��{�O��o\�B/����~�(���B����: ��ao.\C�kf��_@Z��T�\ �͆�v�9��</Sn���k]m��Z�����he�an�P�ݝ�b�Bϱ�[��m�U�H"҆>Xĭ�����̞��>��b��v݋N���������L+-�8���/��:5A��p١w��zj�v1a{J��9H�P�.�}6�/S� ����,��WdM4@�k̇���AG��&'��̞��>��b��v݋N������M}Ĭ���F`���G��k/��m#��}Dq�f����Mڷ��iA'R�	z�#,gB�������&���e�S�[�k]m���E��Y��%�i����w�K��r�]�4�P�l��=5;R�ˊ	18?.���|�T�\ �͆�v�9��Dw\����.m��TDZ��O$mQ��RA��m�q�/��v1a{J�W���]�x}NI0���ԏ�.fOe	m���h������#oM|#9���!�`�(i3N��	�Ȓme":l�nJ�a$�Y ������K�+���w�W���b�0�`
 ֢���뒒���!�`�(i3Ǒ�e}5�,���x!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j&���"�g72O!j���8
�O�@��2��.�g3Z�)V��B�1u:u����<x��u��n�G�A�FC�]s��i�~Fz��Ԥ��C�xi7�E��'Z*)�?�R��nj��P_Q����t�h��W+��W��v1a{J���&Y��V��C�xi7��U��)���Y;e�iK!���d.O.C�U��B��-V���$��b�D ML:���7|)�`�H����Qw�c4~Nr_�mS8<�n�ݚ�Н����D)���Z� ��(HJ�a$�Y dN�<@Iv��nt=:��:5A��p�$�`V1�������S�\zigzA=v)E�g�������(ӈ���m�r����١w��zj�v1a{J��湮��n��>�my$�N��o�/���;�/��@���WdM4@��_�U*�I����~uK7͍��|��W&":�ݚ�Н�K�\7}�W, D�cg�}Ņ��4&Ks�dN�<@Iv��nt=:��:5A��p[�t��#��%��g:���\��Hܞ�E�g�������(ӈ���m�r����;�x'_|~� �S���}me":l�nn��>�my$�N��o�/���;�B�'��a�/������Z� ��(H�I����~uK7͍��|��W&":�ݚ�Н�닓.�`�3BڴQ��J�a$�Y dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3���D)���Z� ��(HJ�a$�Y �C�|J3J��М�Z��N|;^�S;��k]m���r?&��AK��sC宸I))����A�m�(�QNȮ���k/��m#��}Dq�f�9��?xs}�k�����|	�WI�i�<�~�y�j�q�7�AԢ�a\蟴���P`��ʱ�O��W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3�⒍~����v�z`�!�`�(i3���o���F��+=�o$Ô���,��WdM4@��z(�ﳍ�f�_��S�>�!/�_�n�To�[
MQ9�F���"X��[�,�!���D!�`�(i3K�\7}�W,��+G��ܢN��_;���C�|J3J��М�Z�ׄ��e�S�[�k]m���E��Y�W���]�x}NI0���ԏ�.fOe	�b��r�
JB8�^C
��ݚ�Н�[�t��#��l��姹����+�Q�����zk2��|�kڲ��b�Bϱ�[��m�U/|w~S."��b�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J���!<��v�Fr���IbW�P"G�wk�#�_wU|�1Ĵ��ޯi��ŁO�W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3��@�z]��C�x!�H�Z���,ߘ��o���F�������ʂ.m��K�+���w�M�7��<�1�����\�H��/Sg޶��j�}a�cf��"X��[��Q[R�7!�`�(i3�Ɔ ����;ƹ��:i����;qN��	�Ȓ�cЉ�MO`�� \)-�E��%����gr��!�`�(i3���i���w�XU'��
�:qEp�;�P�t�5fĉ>99��A0ok�׹�V���$��b�D ML:�ctj)��>#����,�ǰ?%{B��0B�tw�i�՗[�:X#x^�&����������I �P��M3�G��#'@Nw�z5�0P�ġ��x���u�Y�KG�ξ���I��RhF����u�*��?�d���&�a
�+��8n�TԁC*�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6���n�4��;�jmT�#bs��2[�a��o���H�RtV�^�amf�M '%�줝v)ƍ2���l��k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�amf�M '	��1	�q��eԱ���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��|I����<��}�u�?�d���&��z5�0P�'vr=c�w�N\`�a:-�I�3�BD�O�.r�r+��ސ����U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&GЈH�����b�'Be���0��_�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��lb~*��s��YN
��)e�W�J��H����8�O�5���1tSjv��H�����Ɔ ���Ve��˅�>��{���M�I�h��}�~��l��-/a8!�`�(i3N��	�Ȓ�cЉ�M^�h۾�(�b�'Be�����y�?��}Dq�f������!�`�(i3N��	�Ȓ�cЉ�M�'DV���b�z'hۉ)��d�7�qĉ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�_�Ƭ7~�rG[Pt�����Vx`a"�6�m��gO�J���M���HaU$kX�ڹ��/^�w?�d���&�db�\EX회�h�#5ġ��x���u�Y�KG�ξ���e�J�Pn\�pD��ZOU;��|B���r�����Ɔ �����Vd�;,���3�/�����Y_sĝ���w�R���y�U��\JD:�GI���o�+�=4V��	��yO��aQ'�����f���K�h�y�[ee[V	Q��2�P�?�r�&U���0��PW�%X�9���Ylom;�Ɔ �������4�Ք�R'cf���³5����U��+�Xa�H(�˕�Eo(d��Ylom;�Ɔ �����Vd���ة�蝌b�Bϱ��9��no �گ��h/������B�F~�o3����,�ǰ���9kn��회�h�#5�ޒ�K��6j�"Hs<�?j=Ծ���f���K�h\K�5~�k�좏1Y�����E�����A���@���~$��F��v����{�h�&T�n�2��^�5�^���������EXs70�U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&G�'.�T���Bf����{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^^()��>�����U�._����P�|T����{7�H����8���O�υ���YN
��)e#j�o����B� �b��!�`�(i3���^g�6�x:�m]�c��#���F�H۷`1tSjv�!�`�(i3�T�n��aΪ�;�EIp�r~�h��ݚ�Н���w�w:�!�`�(i36�ZV	�	ҙ���˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�J	���/a���Q=	+�{�*&��q>�<�'���I����� ���JH����8����F)�~����H�V�n8�A�A�y���6���#¯��TG6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3�4br��n��>�my$�N��o�/���;�B�'��a�S���%�����ռt
�AԢ�a\蟟Q��ǺΕR��ӟ-�q�x�~<��w���	�e�<j��.#՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�YN
��)e������p�r~�h��ݚ�Н���w�w:�!�`�(i3%Q�[�J����˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 ��H�����4br��>�=,W�[�?�R��n}�����Hٚ�-����!�`�(i3	�)��&ghRV��R�4br���h�Һ�!�`�(i3��jVѭ@!�`�(i3	�)��&ghRV��RK7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��#}�{��Jw��3��.�g3Zv���� )�W/πs����N�KRK���DV4�ސ���E��'Z*)�?�R��n��h
:h����t�h��W+��W��4br����'�QV[��;_��8W�w��fD�Y%ɫTK���N�KRra?��Ba�Cy}�����:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^���M��2E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����8���d�W�J��H����8�(����T�x�"��XƤ5_�J�	�LÆ���#��p��;�{��!�`�(i32�#���l�
@\ه3
�v�v-}�	mp5���%�+� h�ҩ��wӨj]h���^/e��d�G�.�@��ӯ�2�`<!�`�(i3��jVѭ@!�`�(i3}�1�Ha�E�Rq���my$�N��o�/���;!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���ޡ�m���Y�$�9����~+2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��Wv�A����w�V�"~�ӵ(r7�8� ��$d������`7�tȈ������9P�-�,�AG�<���X饿��!�iv�aQ�Ϧ�M�ኾ���L��r�U���f��/?L���u�D��D1��n������� �k,
"i�̄�ѭ���ɿ�kF��l�l"��l䋬5Kq!�`�(i3!�`�(i3}��[b:��'(K�lc���97�
C�dA��:���f���X�k�J�3���-Q�OP�}.z)y5�[՚1D$Q,�WP����jw8T�1�c�{Wo9�����<��l�Օ��qvdЧ^{�jmWᅫw�5�O�%E#P�;����<��p��b��!���?t��my$�N�����X8�#s�vS�em;����^F�=�_�7V�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��o�.�u:u����<Srƫp��xjzӝ���I(͂��-�����d�tuѼ�!���{��b+}y[�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^>�Q�c6�~nS��\z-+;X���W���b�0�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ����[7Y'��k��F$�kj�L��M����4�	��������A$�P������5d�������y�:Fa�7���W"�P�K¨}�n/�J� &�0D��xjzӝ���I(͂��-�����2��}�����3R�Ƃ�nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����V(MH��ZRR���&���Ɗ3I5=��)Q�]� ���_�hbvk~�#x��Og����1tSjv��wӨj]h��J��sr�lv{��lw	!ݞX�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�ML��M����4�	���P���/��.�g3ZE��g�Hby���=)�Vk����/x �i�{��R�S��>j���T�}ɻY~�y�����[�]9�(b���J��:����}�6�nq����P�U��)���Y;e�iK!���d.B����=1_#u���GT�A�IÙ=�H��'�PD�{y����i�q,?5q��7���9��e���W� �{Z+����"sS<�0�zG�������&G�����$ɔ9Q<ϯ)P<�ܓ�Y�B�'��a���� Ev��\��;�,�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н�|�au�(ZԮ�g��#��ܭ i��Y�{'%sk����w�;F}���V6�!�R/\T&O���GyV�ش�oh��!�`�(i3��=m緒X�X�pF�#}�{��~v� 1��M��%�p@m�ڨ�hծ!�`�(i3��Nh�=f[��8��GM5s�FF���p&1"?�R��n}�����Hٚ�-����!�`�(i3*�9��.���=�⳿P��}Dq�f���.J7h��,?��&�)�
�k\�i��}Dq�f��߆�p�h��{$�������LQ�/8۶&��L�H�W�J��H����8�O�5���1tSjv�!�`�(i3ʬw�S���q9+t�}�ݚ�Н������y����������"��Ra])n#���r�����d�tuѼ�!���{ʬw�S������W�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j �_�ȇLШ��+���Al+�HtB"o
�BP�@Ե5���Wd��%�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6�닓.�`�3�P���F\\���F�`yx�>�+X�M?��y�!�`�(i3�4�	��3|v��Eb�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��lb~*��s�닓.�`�3p��2�H���'T���+8!��?V0D�	�I���_
�u�Y���H�hbvk~�#x�DS�AvF̓@?5�#j�o���&�2����+�+�5���4br������Ľ����Չxv��Օ��qvdЧ^{�j��@�
h����Z>ؼ��XyH�RtV�^q�\E��0�d��+��2VP��Ѣ�ʒN�ċ
�:qEp�;�P�t�5fĉ>99��A0ok�׹�m)��T<�cny��&񮣙�cq@�w�R���y����<�..�4��3�U��`�Р�(�V�'G�+R���o��_�Rv�䩲$��8��I�:Fa�7��X$_V� �6(�X)���7�癆cgQw�c4~Nr_�mS8<�ncp6Dq����Cs�q9+t�}hDJ��3��%�����q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н��xmQ,ۘS���VW��F��+g�ݚ�Н�ʬw�S���<v�cn@�q���uҽfĉ>99��A0ok�����F��O�\E�W��4bX$_V� �6(�X)�ҽ�6jQ����D�X��;���B�9�Q�f�����+� ��*ȑs;��|BX�D�mP�>c��?�B�t�xr�t��b���2�b=���i�WgV}Q
�Waf���� ����6�o8:4�I���c�90B3v�A���('�@�+���3f	aF�o�@OiFA� @D�H*�=bs��2[�a��o���lO	"����q�\E��0Z¥���5.�{_8�Y��=�}�Vݨ�,bxqX��k��^�1��dc�@c�����h��-�����_���`e<�Ia��la��o���lO	"�����2��}��M��V!�D�WaU��,bxqX�HN��R��bP�63Z�t�tH���]*bP�63Z�t����؊O.�x����VǪ =ա�0��L�r:|�O�E/�9��"J j�E��'Z*)�?�R��nj��P_Q����t�h��W+��W�H^��Ƨ�0͜��!?@K�,bxqX�����,�ǰ����E
��sp���m��>#e�6&	  �ιf����ZaL݊���2�"�G�p�Pڹ��/^�w?�d���&��]�o��A����\��]8��	���#�z��%]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M��ŊPTWo9���b��|2\���F�`yx�>�+X�M?��y�!�`�(i3z�
1���;%��v��!�`�(i3��������Z¥���5.�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r���s�Yls��8��GM��-����!�`�(i3z�
1���; ,��rQ�U�^)����ݚ�Н��O)�b�c�!{p85v{��lw	bo N��7�$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��o�.�u:u����<�x���ަ�I��O0Y�6j�"Hs/�n�����E�xc|�+�AR+@|#Z�1�IX0F�MV�ҁGG`5:�����+�^n=\f�5>�.F<!W���t�㮫����"sS<�0�zG�������&G��+�t2�������/��kOT�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*�Va�ir3[�u8���m�~r�D�4�.h=�,\���P�75��iI8�ѐv2�8�n�"X��M�����)m<�3HYʨ�]�_F!�`�(i3��c��qVw���%���RAԢ�a\��?�R�_��sV�����נ2<�i������b��u��r���#�-�p����B��6�<������NM���fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx?�y�g���w�R���yxl+�����o�+��5�s�AEA�W��x�13�K��oNYzZF����9��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7���z�G�	S�uimK������t�r$ɓǃl[�Ƶ�1tSjv� �#0xg�`�I��Wn��>�my$�N��o�/���;����������zՠ�����˦G�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�>��:J�E�<����i"����*ȑs��,:&�^��,Q����-����!�`�(i3R�c4!`��Bf���Q١Ӿ�$���l�K�F���m¡HN��R��bP�63Z�ta�F�������Y���D��3��bt�u�&��F�ߏ��D厺��+�̟�1�8�>r&�G�p�PPS�H�I��I0���ԏ�.fOe	�S�4��=ǚ�-����!�`�(i3Y�)�}��EXs70:���&�����|�b���Fa>t
�:qEp'{w#/ B�d�tu����a{���Bf����{_8�Y��=�}�Vݨ��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍʞ3���h��[��1聦Ά1��<����i"��@#('�cH1��<9Oy��]#�0D�	�I���_
�u�_C�7�2������}0n�V2���]#��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3'����t�Gf��x��9	4��t�f��x���<d3"������-ќv0D�	�I���_
�u�����|�G�p�P��<jV���\�H��/Sg�w��'o�+u�d��D厺��+w���	�e���0��Qܓ'{w#/ B!�`�(i3��7I���|ag��6��+jq����i��gE��[4ҹXH�m�w���i���Z���D�U�2Y��i�p��+˞j��&����Q]� _ό���.�@?d�s�8KFmғO�4}~n���,a�n`5�fK�\w��0]\o�LCd��.ZQ�*�3���g�7s�9���o>��l%i�-}�
�?���B@��������/s9�d�٣��>����C�b!��u�<�`A��_i3i 
�c��]�!����M[��ǢHe�-�c��3E M0�F�T��BZ鎬�����	�7 �#�E �����	(��7�зq8�Ј'���Xw�j�7����w�K�b��2W hbvk~�#x ��M��.ᬵy��"C�����T�\ �͹g}|�H�I��'�!͙��04nԴ�V����U� ���_tE��gVB�3?�J	QT��8&���I�%A?�dL+jq����M~�̀R��n	l��Q;�im��ȍry��	.�n^y���\+��R�4.����P}�=l�q�������g2��Ɏ�#���?�5q{! l��2
L./;�Ly�Af�?ǉ�=�e�MW��Rj�q�wxo�~]�g���[��}��#J*�Rs�08�b(������l__���#���,Wc��I��@�hGq6��nX��U�	vn����R�����_���!�`�(i3#B��F�!�`�(i3!�`�(i3��*�{6��(�w���!�`�(i3Y�"O���j����I~!�`�(i3	�=��G���v�8:ۛ@W:���#���F��n3p_�#2\z��o t�J�PM�Y��G%�&8�,�H*W��u�a�ݚ�Н��^yE⛀B��+ H!�`�(i3ˮF���t�F+������X:��+�i�	��_�V!�`�(i3-��w¹��<d�,��L��#2\z��}�� �с�'(�U�c�&8�,��
�Q!}-[BvGޣkQ�A���ۖ$����nQ�rV,?�����ݚ�Н��V��(��sW��|E�q��w\F��G8T�w�nf�?ǉ�=���S���_�������"�9(���l ��ǣ©���u��4��#�N�X�!�`�(i3�M����iٛ[�Z�Z������s��+qѭ�+g[�</Sn��-�¾L��8�$��`���VF�˷�f�?ǉ�=	s(D��&8�,������	�;�ݚ�Н�4?s����k-����b=�`
 ֢��-�¾L��8�$��`�� ��M�#f�?ǉ�=�ϋ�LΗO�&8�,��@��Y��;�ݚ�Н�*��^�"~H�҂��hWj���H�D���dݮ%*!�`�(i3���_͏��X;p`�����G9L�bW�mT(�l\�6�'����7Z��czZ����N��E�Es!�`�(i3��w]��&��)��>.$5<�`A��_iN��E�Es!�`�(i3)�{� �"�X;p`���2�b=��<�ry^���i�\!�`�(i3�$�~c/v��&EA)<�!�d�<�-�����q$��7�H+�����s��߀������k-�-�����@:[�X�	�J�`Ԡ��`��!�`�(i3��	&�K��2q��'X�qp�c� &��GE<�!�`�(i3�U�s
ƺ�+e;��5&�(�R|�G᭞���Np9�A(jgOR��/�q#a�_�̞��>��3
�v�v-}�	mp,��_А#�<om�����M��2;0��L�r:�9]��j�W>l��? Ah�*h,ChW+x⣗�C��ҷ�㗼�?�S���J8����E^��o۪��5/:�� N
�������?;����IX0F�MV�ҁGG`5:�����+�^n=\f�5>�.F<!W���t�㮫����"sS<�0�zG�������&G��+�t2�������/��kOT�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l����� �'����u��r���#�-�p����B��6�<�������G9L�M�7��<�M�l��S�J*�Rs�08�b(������l__��E� )�&9*�����fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx.F<!W��Y���x�wbk�$ *�������U��RbAvx��բS��\P0RP���50f
V��.ᬵy����� ��g H�8��#eW���Z��1���~!�`�(i3V[B�5�mw�R���y>��yС}������Rr����t70�6�H