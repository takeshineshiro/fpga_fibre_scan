��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�'Y�L(�K�O�{��?f���ʈ�.�֏Pc\֣�I��B���t��|U|�/֚��LT�E�9��h���$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA����q�HS�b"L]$7!����Y�f��a�Z��Vׇӭ��!�`�(i3h��8�|�g"#~j[O\ڀB��+ H!�`�(i3!�`�(i3�f��)<t>���PF�!�`�(i3A�"̙��2�����Vc2�����Vc.|�('��r�dZ��߉�󆭋;2�����VcЁ=�t�!�`�(i3CS�Y%��t[Ed�+֚L��2�����Vc2�����VcϔJCS��G�d<��2�����VcpNR���b,�ҧ�ɟ"Y|fN�:@��翛Sf�\�_�Ճ܇���'o�fqII��*�T�٥��T��|g�S� -E�7*����q��jlw��JF#�dnE��k~xhd����Cr��1��i�Vw�oM �%���bv.�]ֶO�4D6=���i��p�b�G!��Z%�6�ǀg��i��vp�\��M��ڀK�_�rۈX饿��!��o���ݯ_gWgj"���\r��3ة�K�~�'o����֜,ӘkR� �KF
������:��ۜ������;�Ӏ��B[/'g�`	�K4̓������9(���'�Pw��[#M��*�v}���<�LK���i�[-z�g��hs��%�-h���C}�{�c\dnE��k~xnE�HC+��3K�<�s�������5��w�:j�.Ѵ�����T�'�"�ݥQ����2O��'HY-(�3�(M���O|x�Ͱ��Y$��7\F���r��RL�a))�kc�߇���G�/9'�$���'�r{V.� !�zg�Z�$充�pje;��M͝75#S9��%V��"����ʉr���u��w)�Sl���-�ed�~篟|��d���Y��^"� �/Jџ�_�v%�����:��/�|^��D"���b!��k�8���҆�|n����wH�L��Rl[���.���M�ѕ�����aWfL1�Q�j+�B]g������Ⲕ�u��w)�S�3k:�(�-X�7�j���,Ud8J��$�ƶ��Ÿ?%�b8�<�#�1-@��%��Ձ�k�8���҆�|n���)kd&Z0�i&��a�&����?ʳ�W�%"4����*�T������|�OA�
܊��?Y2���3m�!=�y����h�}D�8����8Y�&�\�#�W��a�erp����N�u���u��Uy�PD4KU7B�����<�[0YY���\�4�sP	�b\qB8Y�&�\�@N��B@��2�o n;�q�m���mi=��B�-x=�WD���4B'���S�K��i|ٓ������v9{�$W
?%x�+�� fג�� y�dH�]��/�2�-�]?�B�nI�4q�Qt!��c��<%>ì�oJ5�%,�k�W��T�٥��T�Sҥ��|E�EYZ/� c��(�U����	x]�<���e��8�t��s*ո{�x�G�F�����OwꅂF�-!d6߿��b��'�� |X��M��"�D�u���lٽ�G��k�8���҆�|n����{y�ڋ�jV%[&��\�۱��ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l������ ���yX�ئS��.V&��B֥/~.)��3\�R�F*}�c}��uO�Go@3w��0�c��]W�6�����9&xc闑^����S��������Ǜ�>�xj���+�J��U<o^.K�}�n��&�X&�V�.Ю �{��,��b9���1��]2�?V�Ľ�߉��ə��Q�^�y�zL͊�q��UG�s���q����E©�ʐx�?�'n�^0o�!���!��6�e�:r�"(?�M�_뎱�:L��ҭ�Y�����[�����cJi��2�S�ڬ��M����@qzL͊�q��~���r'�+0�l�R<�q��f�}��h�'f R!�`�(i3c��Et��q���U�ЂDa��(o��0��7�����5	���]���>����C�n��J�
��!�`�(i3c��Et�Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9������>7�,g�YӅ:�v�ј�"��Z鎬�����
��al>���,�۽��E����F��j��\w��0]����jq��Мl�v�ј�"��Z鎬�����	�7 �#�ԬQ���g�z�&����j��\w��0]�o�t���˩��*���]2�y�Z鎬�����	�7 �#�iK�D�b=���>.��j��\w��0]7��u�����a#�fv�ј�"��Z鎬�������(���pl!�6���;b��g��U-�e�,���6+�H�%��ZtV/u9������-��%Mό���.�س���*G��/�p,N�By3��<�]�!��	Ǹ�y85�����3�|#9������q�D���/�p,�]2�y�Z鎬�������(���/��A����Q[R�7�}��C˥�2�6�d�f�����
L'���Xwp�����ʍ�ڑ����E��@IE�U��>��l%i�-�Q�rV�Fg�YӅ:Ԭ����
L'���Xwp����c���i�L�����E��@IE�U����S8�/ #O�)U��֜��3,0=]^	�&|#9����m��
�����\��Fw�]2�y�Z鎬�������(����F�dH�/�R�Ĳ4�������`y�����i�����W��(��"B��$I��w��,c�A�L'Qī�*pY����q�����S�ڬ��MN�ދO�����`y�����i����<)a��/8f�"B��$I��w��,c�A�L'Qī�*pY����q�����S�ڬ��MN�ދO�����`y���C#/<���qg9ۍnJb�
'��(�<��@d�Yt%�)Û4�=w�l��ǐ3����=YN6M�Jv��4�vD�a�ξ���I�2�W� ��iE��G�����(�
t�ژq���U�K͔�����Y�b�Δ;���}�I��w��,>����C��T1�8K��FR��a�z ��(�
t��Y�{'%sAX���	q�KS���K����)��T�\ ��Tǯ�!���\�<�dQ	���qk�ZV"���:��#tCE8�^��㊏')����=.�����b^�'�#9T~�&���#�{�0;�}����\�w�Y��k��ı����V���}���s+���JrC��
��.�z,y�m��P��I��'����cԱn��aМ��IÙ=�H�R����/�R�|_v�:��j��ji���+�z�m_ �e�12Rq�L$�t����C-���&��nX�)AQ������{E���I�$Pb02�O���V���ӕs ��Ӄ�m���VK�4�*�Z�.S����%�z ��y�Κ�9�"�5z���Q��4hz�<Ρ�Jn,���`�rs�i�jf� l��E�4.@�7��y%%��`y����@����gG}O��05GV��#��6�d�٣���N N�S��t�����e6`)K���U�g�q���U�NÍ:��$��fF�:�����,8g5�e`��9����� +��Q]� _ό���.�}�
�?�	�%��6�)r����'���Xw���,D}p$_~R׫��O
'�]�!����w�Հ�b02�O�ّJ8��b9����U_�+X�Ă�L�iۂj2_?.��vœf��yb!��u�<���d1x��r-�T7s�9���o��S8�<�)��'��*�S#^�V]��}R�wX��}�
�?��W� ��iEE���\���n`5�fK�\w��0]b!��uፀ>1J���=������7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���{.[��(��Y�b�΀�e��Ek�Z鎬����t��LJ��{�� ��8D�N����"�,�>E���]�!��	Ǹ�y85�B���0�1���U�<�o���8���/����,Dʝ�o���V��#��6���+�J���q���U��@����gG��@݉_���|�g��s�N���rs�i�kۜ��/�X2�B���s�_��wBW��8���/����,D胬<ċI>%L.�A,���+�J���q���U�h}Nw��農���ߨEc���Δy��Fp����f���,(���B���o��+eQ�s����|#9���b!��u�����Yj<� �1�7s�9���o��S8�<�)��'��*�S#^�V]��}R�wX��}�
�?���	~r��k��by��F�n`5�fK��0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6���2����.�t������:ux����"�,�>E���]�!���X��/64b!��u፵�\�yGL΁�a�n��7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���S���ۍ��9g��?��E����FZ鎬�������(����F�dH�/�R�Ĳ4�������`y���Z��O��<�"��~Ǣ�)�s�ި�b!��u�[��l�,	[�/��87s�9���o>��l%i�-�u��Y'G�~�+yp�l=�������d�٣��v_���Zo��u��Y'G�7s5kL�!�`�(i3�d�٣��v_���Zo��>D��e2���HF3}�
�?��&��>�!�`�(i3�d�٣���N N�S��30���,"�x|ٲ�зq8�Ј'���Xw���,DH�v����ܕz&�8�n`5�fK��0z�cUL���.�1�3�8���/����,D�x ��s��q���nm�n`5�fK�\w��0]b!��u�s�Uo���]H/��d��]�!����w�Հ��}�a��>�A�IS��#�$�~�M�q���U��@����gG5m�E��P����z�7s�9���o>��l%i�-ݓ��E�1�#��d_�E����F�'n�^0o**�ХM
�nGZ��JP�O�?~Gv �@����gG�S���!�`�(i3�b9����U_�+X�Ă�L�i�;#�����v��#;�7���c�t}���#���Q]� _ό���.�}�
�?����S&�r=�������d�٣���N N�S�+w�7�
�p�	%6зq8�Ј'���Xw������LƑ���@�&_E�EYZ/�+V��i|���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�"��B9�
eBZ�tX ��Dsa�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WD�K[�,�ᖠZ�q�PO4�7��V���.g"}�p��q����`U��:
1������Q>ml��B<�D-��I����~u���3rn~{�3�����w���H��(6��W� ��iE��lN���2�0���Q�#<4^��ٝY��e�R��b���T1�8K��Мl��ٝY��e���WDChFb틠���3�;�cM���/���7����*ZV)�J~���L��-aw�n���/�p,�9�+��N�O=�W��Gf��x��9� ��������VW���*	2�f[h�����g.�`�B7d��9�+��Ng�Dp��H�!A+Ǖ�_~�:N�&k@C�Ɨ0z�cUL$8&�{�#�17bN(N���<��D�
�U��r�~�)w�l�-��;��kZ��}.<)a��/8f׾ŞWsuz'���Xw�j�7������on�b�Bϱ��g����EԢ.~���"��h���VG1�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�%A#�@�N�to��h�T� #�3Ł1�q�7��N�6�Q�3u&����J�f���-����R��ݪG�B�	z�M���S�-I�!A(�"#~j[O\�&�����1�sI�Y����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�
t�������t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ�q�� �`>��s��k��^�1��dc�@c�����h��-����'�)�����(9�ϦZ�Be�A�}�	76�&�� Ӗ�t$�)�vx��۽`�$�l,.l&�7s5kL�s�)];I��K�&�a���3Dr+�4���	+��g��=R���>��骾&�2�0���w��_>d�����r�����m:{�!�`�(i3!�`�(i3��!\�'°����ԬQ����lwE��$5���lJ1��j�p�B䁒_[�Ff�?ǉ�=!�`�(i3�#�-�p�m
�ܲ�#���n4s1�U��B��-�ܜr�a���DQ�^�鄃��;��ʁ���MյV~LvA!�`�(i3��w�`L�P�~�9��}Dq�f�}I�6���N�Cٺ��G��Hb� h�ҩ��H����D3w��'��b~*��s�l\�=�]y��d��-��!�"ǉ�t�����J�ϝ�5�v�z�7s5kL�<��r�ŁH�RtV�^CH$�I��*�M/*�3� ���!�`�(i3��\ Nh�gdq�_x�ֺq٫[_�mS8<�n�ݚ�Н��� л�VZ�ڋ���Y�َǤQ�Ї�!�`�(i31���~!�`�(i3����-Jg8�iT��*��C�Y�\�fĉ>99��A0ok�Ra])n#����,����0�|��';��#j�ݚ�Н�VZ�ڋ���Y���GiL�~�fĉ>99��j���GpG�&ց�*�7�|�9��n�7�Y���_j������
C�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^�Jo���jk���%�8�Va�ir{��b�b�*#o�]�ʄ�v�4�?zm�jd7}�� ��M�sv��>���F*a��o���H�RtV�^CH$�I��*�M/*�3� ���!�`�(i3�k��^�1lv0�9l�'����u��r��!�`�(i3��w�`L���ǚ����}Dq�f��߆�p�h�Cd��9s��'}����=��-����!�`�(i3�FW�DVx>74/���RZ�Z]�+����%>�rGO�D mWN՝� s�#�=�U�u�íN=]8k��.ͥ�H�RtV�^pT/�GS�7s5kL������� h�ҩ�9��n�7�Y���_j�����9�x�\M�ݚ�Н��̢k��� :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3����-Jg8�iT��*>������fĉ>99��A0ok��fĉ>99��j���GpG�&ց�*�m*H�	9��n�7�Y���_j����I�����&�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^�Jo���jk���%�8�Va�ir{��b�b�*#o�]�ʄ�v�4�?zm�jd7}�� ��M�sv��>���F*a��o���H�RtV�^CH$�I��*�M/*�3� ���!�`�(i3�k��^�1lv0�9l�'����u��r��!�`�(i3N�-�}q�j�֎����-����!�`�(i3�B&�G���M/*�3��GH�E<5�!�`�(i3CH$�I��*�M/*�3� ���!�`�(i3�	��x��ݚ�Н�9��n�7�Y���_j������
C�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEpj�E}4ظ�N�Cٺ��������� h�ҩ��H����lv0�9l�'����u��r��!�`�(i3��w�`L�ķ@���k>��}Dq�f�HN��R��bP�63Z�tHN��R��F F�E̠(*�O�q�)����CH$�I��*�M/*�3��GH�E<5�!�`�(i3����,����0�|�_�mS8<�n�ݚ�Н�-��)'�>���F*a��o���H�RtV�^CH$�I��*�M/*�3��q�t	<!�`�(i3��\ Nh'{w#/ B!�`�(i3��S����=����h�[� �c��!�`�(i3��Ě�����}Dq�f��k��^�1���+1��*Hx�g���-����!�`�(i3Y�5�n�����_�������&G!�`�(i3VZ�ڋ���Y���GiL�~�
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W���{��s�J��ݚ�Н�����-Jg8�iT��*���a���݄�倮(���������d9=���u��r��;�jmT�#�0M�Ŷ�Eʨ�`N/������&G!�`�(i3-��)'�>���F*a��o���H�RtV�^!�`�(i3��w�`L�P�~�9��}Dq�f�՝� s�#t��ۻz�˾ �����]&�U��f�!�`�(i3<�6�Q=�hNNR!���	�-�ud��X縤�q
˾�'v����UrSuͫh�<���D��ܒT���.�[M���r����!�`�(i3�(�d���Հ�ˤ�䁔�`i�����tZ>P��]�{iK���	����;� �GE@��!�`�(i3VZ�ڋ���Y��ˇ*�h��!�`�(i3���F��O��ݚ�Н��̢k����0M�Ŷ斗���%�������&G!�`�(i33~��d�Mkٴ�$a�DkW�����JӉ��;4e!�`�(i3���ܚ��@��f�\%�~��\��8!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����V(pyL0DMlE'�! CH$�I��*�M/*�3��7ݽ��!�`�(i3}�	76�&�|��3��׹��ܜr�a1r8���I����ht��ܜ�[�^���H> �D�9�{*�,6����Z9��J����*��m4�b �	H!
�I�N��M6f��,�,&�J�����7�y��ħ���n��$z.��X� 2!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i33��0�����+1�;�.��1���,:&�����9�Ԇ��|Z�.!�`�(i3!�`�(i3v4{����U�ɶ)Z�_v(��ڥ����Ⱦ��,Յ�1���~!�`�(i3?Q�@X>#�-aw�n�W�^�|��p�@OM.Ir�H����2��b�Bϱ��>1J���� ��0� 1���~!�`�(i3?Q�@X>#�""Q���S=�r?z�3� �mKgN�쁘o	�V�6�J�J KB�~�.$d�I�vNR[��j��d��\\N�2߄��`c�N엁�7���R��4�{$�^&��AՉ������b�Y>�fWj�t�[LY�ЈɄu����0��|͖Dzd�=�/�t��Ǽ�d%���P�.�5k��~��/6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G'9�и��{4hz�<Ρa�E�Rq���my$�N��o�/���;�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#&�|Ξ쭧S{#�lܵ�p���S��íN=]n�|�-3�lv0�9l���ў�L��X� 2���t��Һ'��b�%���!j�l��XulMd�[���}��M�?L}�7x{^4��*m!�`�(i3�����V?��	����pॻ}����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍٽt� $�N�����"���Q�������t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ��W�3�-6�n��j&b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����Zj���
���+1�;�.��1��!*��*8��!�qg�L�[\�"��-����;�jmT�#�[�#��w� ��Ք��ݚ�Н�U��p��PrΌ^pG2��$�)�vx�;�U4�IgWaU �IH�RtV�^>�Q�c6�J�
�Mɏ����V?��Ht�!
�:qEp'{w#/ B�d�tuљ�FdG@/X��-�����+Ut���$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�qb�V�_2��Z���}��C˥�ɗ�iL�G��IX0F�MV�ҁGG%4vkz����`���φ��<�6����N4�,�7����r$ɓǃl[�Ƶ�1tSjv��[�	���d�~{��)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���]���`T����+1�;�.��1�](g���������lҡ"#�k�d�8��k�SA/��M����,�,&�����ᇱ�@�=%��d��-��!g��J�s��z�
1���;#o�]�ʄ�v�4�?zm�L�[\�"s)l໶�,3��0���3i��U��N��M6f��,�,&��$��!'Q5/�dI{��XW���!�`�(i3+��Fe���5��o*4�"ǉ�t�0/0`9N1&�2����1tSjv���������5)��Z^�h��N�M�ob�H���T�ì��������R3Y@T���אQ�B�<}׼����!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3U`�Ȝ�W�iy��*)ci���{2�k��^�1�3i��U��8����q �H�%��ZtV1{,�m���B� �b�Ћ����$�~�+yp�l���d�L������.��U)�~[��Q,��:5A��p��jVѭ@�mJ�0�6������$�~�+yp�l�#QSU:�����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�+	=H�ลGH!aߗ��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���
�x^�LRXN+EWE� �����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcZ�)���,I�$�*�����t�T��?E-h��`f���sd�G}%����3f۪�G�Q���x�\���F�`yx�>�+X�M?��yЕd�tuѽ3y��s��>H�,b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-����>�Q�c6��=�ڹ&��nF���<�W�.�P�	��
�Q�}Ql4�u��;	ȕ?�'����u��r��>�Q�c6��=�ڹ&XC�K�7(��gY6!�K������B�̢k���`&c�'N�jLm�<o��M?��y�!�`�(i37�UyR�j����^7��œсW��e�p�x��;b�-�2��|$*g!<�A�IS��03�� <I�����&G�����$ZtgQ�9OZ�s:�8��z�Ȓ��\:9�C�s�4���%>�rG�@�	����$f��_Ub���uQL+��φ��<�6�l�x8��-a=F�!#�&��>�quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\70C.�>��V�m^݆��xjzӝ���I(͂��-����J>zߋ��>ַ�����ƍ2���l�����g�Z��3��a���!@�f")u��r��}I�6���N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s��m���>G��Hb� h�ҩΞ �@[������4Yz����|e"���F��O��|#HK�� ��5%q���f�e�x��w����֯���,mk��L��a�	�Z���ވ��*I���b�Bϱ��>1J���� ��0� 1tSjv��l�de����O|���/��kOT$f��_Ub��7��G_���;�P�t�5�׹���8�2W6�[�6���"����)W[�ۺ�E�`�4�l�T�܆rl���CLmk����������B�s�Uo����~c��0���IX0F�MV�ҁGG%4vkz����`���φ��<�6�`&c�'N�j��v�����r$ɓǃl[�Ƶ�1tSjv�œ&|�9�n��~��4�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b�Ѐ�(���0���;	ȕ?�q9+t�}�|#HK�� ��5%q���f�e�!\���k���%�8�gVdxQ,#�%+V��t�v��ONH!�`�(i3s�Uo���ַ������?D�8����Ě����E�i�m}6O�D mWN��ܐ�}ĚȜ��Y���ۉ��K�A�a�ܥ��(J]֞��_�TYh�p��_����3Y����P-r�uh����s�Uo���P�<�^�s�IX0F�MV�ҁGG%4vkz����`���φ��<�6�`&c�'N�j8D�r^�Hd���"sS<�0�zG�������&G��(���0�l{�]&"(�q9+t�}����@|����^a�nu4Bޗ��jw�	�����*y}e�����ӽC�H�CW���|e"�K�,ǆ�`�íN=]b~*��s�h3pX���Ь�J������pك �%�K��^/p#��I2�8��[�@���=aS�H��ݚ�Н�`&c�'N�j���$�a���NM���$f��_Ub��7��G_���;�P�t�5�׹����忔8l{�]&"(��0�"�˲yQڥ�#�Gւ�Ѓ0�ߔ�;�&���b����~�]��/�\����P �"ƾ��gx�׈�xIY��8>h�|�Ȝ��quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7lk�p�+N᢯��0�8D�r^�Hd���"sS<�0�zG�������&G��೹�C�A�IS��[;\v�a��ƍ2���l�����g�Z��3��a���!@�f")u��r��Y��8>h�|�Ȝ���q9+t�}�|#HK�� ��5%q���f�e�!\���x�sl��Va�ir&�����2q(���27:�������&2��OY�J�M����!�`�(i3�Uʮ�V(Y�t���1�g״$(�>g�fĉ>99��A0ok�����F��O�\E�W��4b�⾰��bK���żh��e� S�p���k��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�sݸ�/�gxjzӝ���I(͂��-������!�����ִ���	ɩ���@|����^a�nu4Bޗ��jw�	���|#HK�� ��5%q���f�e�x��w����֯���,mk��L�������&G����l��>J��Ëf���:�I����Q؃�L�/�Ѿf��6�$VV���ݚ�Н�ٮOS���pޣHV�v&
1����nX��-/a8!�`�(i35i�a�vb�^օ?D^��՝� s�#���k$ '9�и��{.��_+��y�և@>������$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�6�~�q�
4������; i�V�JD�IX0F�MV�ҁGG%4vkz����`���φ��<�6�c��:� �����"sS<�0�zG�������&GU�z���K� |�>��̢k���F�KD�Vr[/}>5��0�B� �b���H�������3rnu�j�fK������&G����l��w�|l�>P"G�wk���zܳX�P��%�©p��;�{��!�`�(i3u�st����'�PD��	��x��ݚ�Н�9O�m96�o9i�!>������$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxyk���]{�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�{�ը7�<P�qb`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �,�E�ϣ%�t�/7��[��IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��y�H������N����n��>�my$�N��o�/���;WJ�Vп;3�����I����~u/��kOT=�40]���8�C�Ћu�a�E�Rq���my$�N��o�/���;#&WJ�z�6�2�^�?�/��kOT*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t��[���}��M�?L}�7�����&G�0�9&،�Zg�x��J�a$�Y �c��~����}Dq�f�u��y\G��&N"3A�NO�]���
 v�n�t{�k����l��e޸XhZ$�2p[_��bݯ�Z ���vت��ݚ�Н���m15sV��#��6�g�.�n;c`3jYYf���%>�rGO�D mWN��Ě����ڻC�i�φ��<�6�9Ϲ{M�9���	��9e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!$W�j v�H��r�22�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc&��!��Q�a!7g���t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��y�P#+_]ݱ�t�UW���.E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t�	���QC�꠼*d�m�d��-��!|�|�����@��pr��4N�J�ף�<Jq�Z9�`u0�F��a�Va�ir�À���<��aEG���B� �b�ПB�'��a�e���F�&Q@d�ݖξ(��D�̢k���
�I�8����q �H�%��ZtV1{,�m�ښ�-����P#+_]ݱ�t�UW���.2h+�qGR�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b׏����e���F�&�c��fly�dCn:�l�U��)���Y;e�iK!���d.��$�Qu�G���z銨���`!'���Xw�j�7����w�K��ݑ�][H5���8�R�wX��d=��¾ȼ\���F�`yx�>�+X�M?��y��M;<QA�"�pM�00_��nF���<�W�.�P�	��
�Q�}�1�:v�!�ӛu.�A�e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�m���>#o�]�ʄ�M��,����q���f�e�x��w����֯���,mk��L��q���3�tޙp���/�dI{�n�|�-3�A���|���d��-��!�"ǉ�t���S`5�㬌�$Q� �H�RtV�^�\!�U�o�uр�_�mS8<�n�ݚ�Н��B*�0��If�<��}��ŁAm�̞��>����� +�z���a���Nq~o@��b+}y[!�`�(i3�g����E�r)1;�Os�rs�i� S�xSVe�f���,@4!F�0�pD8��a�{�
�:qEp'{w#/ BoU�� @k��m�pURƩc��~����}Dq�f�"�a�BOPj�+*7u`��]�!��	Ǹ�y85��X��I�ՠHu��0 H��B�%V���:5A��p$f��_Ub�F�S�1 �T+���f��,�,&��`�2,�!���������d9=���u��r��Jo���j�"Iե��G��Hb� h�ҩ���YeԿf��&-Q��������M�7��<��am��	t�O8��4a(􆿳���ʮ�����|e"�c ��4�-+��.���!���c�A�L'�ɻ�}?s��{�2V���ś���k��	��x��ݚ�Н��B*�0��IT�q��]7�Zg�x����}Dq�f�"�a�BOPj�+*7u`��]�!��	Ǹ�y85��X��I�ՠHu��0 H��B�%V���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx���$4gozq<����Re��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!$W�j v�'���H}�@v���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h;�ƽ�/����zN�S���t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��y�P#+_]ݱ�m�
���nGW�:!�E�/��kOT*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t�	���QC�꠼*d�m�d��-��!|�|�����@��pr��4N�J�ף�<Jq�Z9�`u0�F��a�Va�ir�À���<��aEG���B� �b�ПB�'��a���{y�mV8��0��1�"�"��K�w(T"c!s��̢k���
�I�8����q �H�%��ZtV1{,�m�ښ�-����P#+_]ݱ�m�
���nGW�:!�EҰ�WDChFb�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b׏������{y�mV8�	՚�^��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������]މ�;�Gۍq��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!@+�ϕ���q��B�`�J�ɉ�z=� ���ɡgJ��E&(p�
�Eu�J�?Ig�(��9��ᩃ	tN�\c�-2���S&ϊ�;ѩ�E��p��u��.t�=EpH��j��A�0: ��q����%	�3)���C*4��]���
@�i��g�?�d���&�V��o5]�:�b��t.�C��6�o8:4ښ�*jl���C>��ӚH�RtV�^����Y�z0=�_���{_8�Y��=�}�Vݨ��}Dq�f��R'cf��>��YfG��-}RY
xǍ�J�r��ps��u1,����Uh1�[��(��;�jmT�#PB��/���߰�$|�Pu��r��;�jmT�#��	�DůI�߷�c/��-����!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H��Ⱥ�Q���'g`$�YD ��� ��?D�8�鉅�%>�rGO�D mWN՝� s�#���k$ �H����ڻ�+���i��ċ�!1tSjv�!�`�(i3
/���p\"�!˥���KS����<;�$��\|����=�'�^�����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��?�JY�)�,�Ջ ��C$�)�vxZ`�b�0P!6j�"Hsކl9�p��e޸XhZ]<�����	��TtU��
g1�MVjg[؎��&���.ԥZs33� �=X����\�5�O�%E#Pʲ��U�4Y9��?�s 90� �p/�ϸ<��F���m¡�`��&0�yl�q�����U��)��~0&ۅN,d@�QMA���8-|�D�7��aM*:�b��t�l��p�xB�my$�N��o�/���;�SENan&�� ���� �KS���*�oF���cԱn�+|�[Xs�g��������:=�)��S�2�]�Q$iP����p��ݚ�Н�X19�-.|}�$V���<M�~�K������&G!�`�(i3SݳD��zJe޸XhZ��-����28��m)[�Z(V�eQ״$(�>g�!�`�(i3���F��O��ݚ�Н���jVѭ@!�`�(i3i}B2>�~ə������'����u��r��!�`�(i3����Y̀�3#O�2�B���s�����X�X���`��,n��뾦�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�fF�5.]���E�i�m}6߸��S�Ȍ��9�ڮW;��|Bΐߧ �l�}!�#�b�$2j�K_ryQ�j6�S�z�����F�t�ϛ�c�.[K��mZ�'����Z�G�a}C��B�No
/���p�U�.��k��~��/6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r��;�ƽ�/��e޸XhZ����xO<�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H����D3w��'��b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���܌��!���uxrBZ@2`u0�F��ay�z�v�À����@���l��[���}��M�?L}�7;Ȼs���ݚ�Н��T1�8K��}!�#�b:��c&<:�b��t�����W��k��^�1��[��o}��MX�w����D����K�f�1tSjv�K��ft��;�cM���/.�,/j��O�`�mp8V��%�TgR'��}Dq�f��5ߧE4��mJ�0�6�$f��_Ub���uQL+��φ��<�6�
/���p�U�.��eWo�A2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܺ����ܟgx�/.ؘ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������c����}�I��}ܚփ�c���A�N��'���#����x��_�ΙB5��~�6�o8:4ښ�*jl���d=��¾ȼ��C7}n���R�E�g�������(ӈ���m�r�����i7N�_�Ar��� ��w�K��ݑ�][H�#Sv�Dr3�'g`$�YO\����*A&-�Ri�)��S�2�]�Q$i��a��ݚ�Н�����SP��'�K �_�mS8<�n�ݚ�Н� b��tY�0�����V	���Ċ��NM����Ra])n#���r������C7}n���R����c�Q0��b+}y[���%>�rGO�D mWNHN��R��bP�63Z�tfF�5.]��aT��3G�IX0F�M���3�#<�W�'�B��"Iե�䛑��e���kn%���-j����O�ct���|��U��'"!�U��)���Y;e�iK!���d.���+�^n=\f�5>�� U�c�pl�Ф�T���r$ɓǃl[�Ƶ�1tSjv��m��
��>W�~���%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�m���>#o�]�ʄ�M��,����q���f�e�x��w����֯���,mk��L��q���3�tޙp���/�dI{�n�|�-3��e��2
-�XC�������,:&Ȍ�g�F��6�2d�I����ݚ�Н��W� ��iE��h�{:m�vW(�����C�Y�\�T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH�H�߳Mk��{	�*Nx����O�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�]~j�wҍ���]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�`c�N여��;�Ӏ�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0�]y�Q�'��3#2Ex��D{��#!��׏��Z�׽i+�ȕW��L
��^օ?D^��MQ���0f�Ϡ�����b+}y[MQ���0�-��h���i!��6j�"Hs^�Z�cY�Z��~`a�K��j��A왏3#2Ex��D{��F���ˏ��Z��C#/<���q6 fd�i��sM}�!>m�Z9a\�-eO��v��èb|5�;l������Q"}Hi��v����o�A�,�
=���f�,�k]�c�jd�L�N��Ưb75���J>n�	G0��t�UW���.@�n������O%��}|�[]?=���N���9����v���V������yآ�D�����尠"������d�bv�h�C��p�@OM.Ir�m���>#o�]�ʄ�M��,����q���f�e�j�5˺����D���.���z�<,�\δ!�}�fb���l!c�ڀAԢ�a\�2}$#h6�ćm'_��Mw#�vzR5�<���X��O���r����!�`�(i3�>d�g�KR���8��h�	�O�zφ��<�6�@a� ��fFMqlgd=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^MQ���0�-��h��ƍ2���l��k��^�1��dc�@c�����h��-����<�6�Q=�y'��BS�6n��e�<y�������H ^muN��A`	`#&�Z��1�O?rof�B�
�о�J<������j��H�߶:�3���.�BU�h����;��#�a�Ą�����kO�d��-��!$�)�vx�;�U4�I�';��#j�ݚ�Н���f�,�k]Cw�Hm��/��kOT�Ra])n#�ґ`�g�y z�P��	���QC�íN=]b~*��s��ݚ�Н����a�so!�}�fb���l!c�ڀAԢ�a\�2}$#h6�ćm'_��Mw#�vzR5�<��KɸǑ��)��#���?{����;�.����^����>=���#u��r���#�-�p�G�6�!~�n��뾦�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j�@�f�smy=$o��ɝ1��,Ƌ��6j�"Hs#�{'�?~o_���B䁒_[�FquA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7�p���"Fi���*	\���F�`yx�>�+X�M?��y��#�-�p�%��a�����b+}y[�k��^�1��dc�@c�����h��-������#�a�Ą/�dI{�b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����-�����#�-�p�%��a����"��ӌ�rHN��R��bP�63Z�t��m�5h1���g�F��6&�U��f�!�`�(i3b�6��R%��v�ډ��%>�rGO�D mWN��Ě���aT��3G�IX0F�MY�J+�WTI�;}it�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc4�`�(H��L����M�,!hޖ�A$�P������5d��n4s1�U��B��-_S���\��uW������r$ɓǃl[�Ƶ�1tSjv�t�R!ME�'�^��������@|����^a�nu4Bޗ��jw�	���|#HK���4Y{]$�AՁ_�mS8<�n�ݚ�Н���Q7lY��)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b����A�ձ^�Qb�Upq���!���_2��VU(��z�j�Aa�R�