��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�յ�'�)���Ҷt�*^��I�.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo�����(����5���&<˴m�mPۑ��X��]P*m����)O��Ξ4�"�\�� ���K�O�{�����8�\�3��>M[c\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�(����5���&<˴m�mPۑ��X��]P*mQg�@zh�S҆�|n����Շ_ Q -���W}�+��X��J�Й�m����u�����w`q�tc�ؑ��g�=Iĩ�m��d�7�Q����.P2:}��>�,�_'�hQr�k@Q��j��C�뫰v]uR����Pl����N�Er��xXc)O�%���ʅ�$n��RL�a)=�y�~ ���G�/9��i�:��^��I��X�7C��H���j�v�?�*�u��q[o��>�`u^9�렕4��S��$[��������\�4�sP	�b\qB��������"^Y怄�GW���և~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��E{�V���/��aG�k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"�~�#�B7#�̔"v��ƒ)?˳ea�8���?_�5/!�"��3g�ݜ��q�©���d��P��}()pxt4���J4xʆ�ĲW��,)B�|aڧ������'Sea�8���`<4}��(����5�2���[@%����nEA�i�+���NؙbG�Jlf)@̲#�G%�&0ĳ]o��in�m��+ r���7����^�L[ b�����,\ަ�It�k\,آ(��XK��(ڷ|��'�u�'n�^0o��~+�ݗ����Kp&�@���k��l0��F��jT�����N��3w:��O%��<������4];ˍH�F�� g���t�&_���9��E����F�'n�^0o��ҕƦn+0�l�R<�q��f�}��?��[�<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����(��eظ��7�
BcyMu򔲊'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5��6��	���`y����ꢤ�Og�?�#B,�Ң�{l�f|�m�jp=�>��o�
�v�ξ����LUG���>��Oޏ��F˯�+)�"j���b7|#9���{k�h�++k&v�Iz7G#+�ǚ'b�t	�U���C��O]r�<Uee�,��3�L���&Ã�M�R�^Ƒ�Өg��U-�eaԗ5��C�6�ǌ�lA�1�:�Ω�յ�'�)���Ҷt��Ah$��>���67�a��c���}��D���(��z�j�)�q��1�:�Ω�յ�'�)���Ҷt�9&xc闑^hY����r�;*�}Ւ�~ܔp�l
d�o�R�N:��,��g�7�s<��MR�������c�A�L'��!�a��5�%]���a(􆿳��?ƾ��s�h�
!7<���������	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�/ #O�)R�^Ƒ�Өg��U-�ez�r�6��DP֞ >�@N����;*�}Ւ�~ܔp�l
d�R�.��On��M��������4����/����DP֞ �+DB4O�;*�}Ւ�~ܔp�l
d�R�.��On��M��������4����/����DP֞ T{o$�m�4|*uN�wHZr��AR1<]Q�I����踫g(�r��!9nV�[}�@��LJ�W��7/��T:���V��Ϧ�p��!K��tf��
_�n�@/%{�;����f�kN�ı��XK��(ړ�8ݻ<�_���,D�i?��Ǚj��4oWpH7���
I@1�ؠ&���Z02��`�z��4�+|'yG`ݜk�@����gG��������&�K̶*|*uN�wHZr��AR1<]Q�I����踫g(�r��!9nV�[}�@��L�ȓ�iӚ/�����&��)����!��`,9�H�W��`�z��4�+|'AB�c�0����Z��q�\E��0Yeώ�$ʈ̷_��yC��S8�dQm��n�R�W�6?��D��~u��v�9��(�H�`��{-� �y��'���Xw�j�7��XA��N���I���X�������/z*q+6j�"Hs0�4	�!]�/)���w��� e�V���<�G]���³5����XK��(��s�Ӻ���?�d���&�	���DLC�Q�K� ID�c=p����������js[��J��:����a�0�I�̡Q�1�����F�+g+�'���Xw�j�7���W�6?��ycP��$m6N8]�؊�, ���q3HL�1p/-��� r����XK��(ڿ�[���7[��}�.���v�9�ʜ���,�ǰ�f,�Ob��^g�MPǟ$y6:[�ҝ��_'�p�MŃ�,��)ǆ���B(��@PM�5�O�%E#Pl�i�<�9��ݠ�.���?r$��Z鎬�������(���kO��u�}���	�f��/�Pqh.X��#�W��'�)�Բcf�b$j�p�t�v��I�`2ڻ�Ϊ���&3�{�H���~��w�R���y�\��ǼPLɌ�Z��E��3?�d���&���Ȩ[�0�X��(!HX��oȺf��[��a��_?�d���&��r�2����^1����հ v�	�أͽgF"?�['����?���F����H�V�7�}�!���Lr}��U�o��_�Rv�䩲$���dS@Ɵ�oC>��ӚH�RtV�^xjzӝ���I(͂��-����!�`�(i3��,� �݂��\���/dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�B� �b��!�`�(i3y�}�6f&rG��Hb� h�ҩ��wӨj]h�,?��ri0������q�+�TM`�Os3�����:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;��mךBo�N���
H=V��	��y�\����2�-՝-xC�;��|B�&�cD+�OW��9�.�8{���@^�4���z�k��q��־�W+��W�e�v��ҵl+�TM`�OaT��3G?�d���&�U(��t*H����]��� n`Ip�\{ف(�7���<��Y���XK��(ړ�8ݻ<�_;��|B
y�3~;�>o崭�kvWދ�qc:`$�P.eE������v�h�g��U-�e a⣃_B7�}�!���*��]o{��#ɱ�|w�{P^K���t`x;�}Dq�f�#l~+� ��IKc;����ef���z�?Y[#g��}�	76�&�;��|B4<d��
~aT��3G?�d���&�[�I�WꐊO�A4ZY�j(&
M�K;��%YM�	�v�3��!9nV܁�8y�Ɋ�W�w��fD��3�l�=�g��4� �㎿���o��A�q�m�,���P�7� �g��U-�e a⣃_B7�}�!��+��%�k<ꬺ��1����t��PЉ�Bk ���E�i�m}66j�"Hs)H��4)�>�|NU�jRV��	��y~��52�0�C(�M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��(J]֞����*/�|�'ɬ���`����
��f%���ܴ�>��}l�$\�U��v�Ɔg��;��}Z�
d~~������ ���tn�u�"LT߫�%��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��VH�nEsu$�D��=�U�p�[����������y��=��!�`�(i3߼��� ��Z$�j]x�7c�oW��mJ�lR�!�`�(i3F��|�'�&퇖+rv�a�L���$ɀJ�ߒ��@���?6�!�>��2%��0n��1�c\ t ����_��V�0]p4s�m.Xry�~�fh����爮��J��ڝr�F`�k��m6[��-�b�+�