��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�L'jf-�6U�P�H�q}^������=���u�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k��O��ڴ���WЋ��I�?g�f�ja1�n�[�ެT�Z¤��I^��?�;��XC*^��I���b1Ø^���#K���lӧIA�a�V��R�}9����3�c��J�'�دv)h�V~�$v�p��"}�v\-8�������>�`)���a��rl�ʩ{�Bf��� ��|4�VDG+�������X".��>��'��E����F�Rm�I�|^�Q�;(1Z �bRw�����IL�+�{Dr[��	�� '�T�������3�f�_��ic�n�QX�v����<.���+��T��/o��إ�8p	�rh5��tE�ӻ���Z=%�-ǋ 4�i� ���������	x]�V�����v����,B���_ġ��M�S�O1��*F=ॵ�h��!`Þ3�����c���.�6X�,4�?n5���AQ� ;-]6�*20��K�X��=o����"���	x]̍�9��H��@N?�qt�-U��S���D	��e#�'���'�A�n���Bu����\�4�sƐ�hd	���Z�<uoѼ�=nq���i}3�L����­��+X�0�w�Gu������	��wˏ����J�2j���_��J��RL�a)'r�Ӟh� �������JܠR)1���;$�� ֹY���8hjY탌�S[W���9��1WA"SӠ�|&�q�!h���噞� x�����Kr4��n�:��e]މ�;���J�	�هU7S�>
��W�Qx�ـ� {�����G��D��;B&�� �=�?��"�Tp!!v*!��1�����f��{0��d# c��(�U����	x]�fX�eϝ(�&Vi���ܩ[߹f>N�u8t������kk��������yȝ�No��>���:E[Kڱ�cTm�Q�����<D���Yl�2���[db���"�p�����J����R�"+���Ŝ�g���
� �AH�W���,v����,B�_�>��\�A�D�S�O1����l�n�Zl���H��6֛Q��RP���敿���|q.;�aE$ /j��sZ19(�?Z��pV�����U-�P�?��ԭ� � �n^�*���j�Ƿ�:h�(n c��(�U����	x]�<���e���٬���f��S���D	����,R�/�G�m!7�X��@$W�ػ��Y�׍�C�	9�/{�ڌ%|w�u�]bu̎}�Zq��Ь��dy�D��3	�53�'6��
�U��p騥m�!=�y����h�}�N�5�%���3�3� ֪-H��U�)��NT[�����=��A|����n���g��k�8���҆�|n����0ӵ�q�TGWXR�� �*xf�+���B�x�
�b+S�������\�4�s��{��]Qǯ������(2�SnFUR�.�;�~�MUs �9�N��U*��$1Xf_q[o��>�`u^9�렕4��S��$[��������\�4�s|��Z�w�N	:.���nњ�@I�y���޷����7C��Hc)𡔚I<Y�@�Nq"Jc�l�!H���uS �����g�Y!#v��v�0gSx̏7�ɍb�e��}vh�xC��6֯�x9���z�{AN��L��xScKE#���,��n��zWi@�!����,x�}vh�xC�}��C�p �Q8�m���8��!�3".t�|6
~����0_�r�O��C��0������m�Q 0��]�������n�u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L�S5H�j.F�k�5��Y��{��/Ƽ���\�4�sƐ�hd	�ѕy$h��ݔf5*`]�|$ɋ��c�~�MUs c�+պNE��#Y��#p��'��������S�����:�֣I���Y/��S"�:����:�wl B����/��;��|B�6L����k�y.�)$����\�4�smg�:�TZz�xy�V�
7w��C�QQ�mqx�F�~�MUs �.Eٓ�9PHvE�	��5j�rO�r�O��C��0���A�w"�mߍu�M9����)�&�3ԫ�쏩7C��H�Zx��%Q��q�\u7i;���35wnq�M�4���d|1l%�<D��8�Ӂ��mw|���^��Bc���pQ�U�.��3�����^"��텿6>��PD$i��^�aB~�q�M�4V�ZHSB�k�� �9m�!=�y����h�}D�8����0�.�	�Z*E��n�.n��vs!��~�MUs z�\v�Ζ�oK䝗�EJ�{,;!Zќ���ǣ�"n8$[RX'W�=������Hw�Q�[K�1a���t~k���a� ����\q�r�"Q'MH�kX���7}p��a~r�O��C��0��`�R&.1���L.��+�ד�4B"��u���;��l)P�u��]�@	@�Xn��r�O��C��0��0RC��L����H7�^��k���D���H��~�7C��HZ�[�0�7٢z|Mߘ����g�/@�G��P��\�4�s���rH
>TT	q��$�2�����b��ǾI}`�~�MUs �?oQ�%'�s����o���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�ĲW��,)B�|aڧ������'SR����.�}|��ι%9T��7���S5H�j.F�YZY0@ìO6�Pr"?D2BC��5��Yk"1/���%	v3�.�z,yI�k��S�����ˉ�1�:�Ω�=A���>�L'jf-�6U�P�H�q}^������[ b�����,\ަ�It�k\,آ(&l������g����=l0��F��jT�����N��2�F�PǙ#Y\��?�l~�Uf���}��\�v�T?�7G|`�UxHj,��|��	�"�,�>E����\�v�X�zgq����2��̪U��֜��3"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3JHn��z�_c)���8���bg�1�Z���=�������b9����,����d���z���ߘ�)�I��<
DN�l0��F��j�q	k���A���������]c���H������i�=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3���D	��U�l>o��|�,+$\�M���j��"n+0�l�R<�q��f�}��Gظ0����!�`�(i3��|g�Y�'���Xw�f�VHF��Q�#<4^��E����F��j��\w��0]�\�LtF�!�`�(i3N�By3��<�]�!����M[��Ǣ�<��>��%@��4��c��Et�Y�{'%s�[�&B�踫g(�r� k�|6�8�3 �;]�F˯�+)�"j���b7|#9����nސ��3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��Vx�%L��W��_�ړ8���/����R�Jm���S�����*���j�Ƿ�:h�(n�_cn��\N�2߄�2W���R0L�>��0�]2�y�Z鎬�������(���_U)�<�&#R�^Ƒ����"X��[s�o0�` s�"��=�6��w������
L'���Xw s4S�'�i��`�z6/������,���eFz����zf�U����z~��6��	�\�HP@�a%=dϖ�i�@O�x�7���q�©��'w��
�fʖG�œ����s��3�m F���9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8���	�~�����F��mF�!؂�����%�}< V�5��D�of�7���A3�(N��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L�P7koеI͢'�����t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s�h�v��T�v��1���6��	���`y�����������T:���V��2�k��in>����׌7<���������	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8��L���NQى�m)k#֫��/f��Ԝ�]����n�4�{lGD�V�B��иܖ��A�.u�r����.�p�m~|��8yL2�����ތ�1�"5� �S�n���&&�F˯�+)�Pg�����R�^Ƒ���P4ǲ �n�/?S�+���LQ��b9�����:�{��ߘ�)�IF��M�����%��/q|k��԰�/"��nH�W��b9����2�u|�Ǚ#Y\��?�l~�U����ۤ�
KlG&�P���ei*������5���􋲜`�m	H��|����OxtX+�Y��M��ҹf�f3'\l�'$9��`�[�*!-R�^Ƒ����"X��[�d�a�4$�b!��u��<��>�ڃ}0�z��D�of�7���A3�(N��㎏qló��@d���/��=��K�R�hE!3�͸@����gG�DI߃��S�*;qܕ�'�e��`�)�	�%{�;����f�kN�ı&l����[}�@��L}�
�?�G.�:��@B!�`�(i3��P>Z���`�m	H����5b11��m��0�]cJȷW+`�x�o%t���,V=ri�{���иܖ��E����B���qEـw�"�Hߢ�]�C�K��ƃ
ᾆ�x�T�\ ��y�.�`L��DtD�z�����0��V�6IWJE����g�%�H?�Q�q��ʃ���_����,D�푧)��k��4j�^oP��a�I�pukZ��@`� Ei�lmZYQ~�H:�����|!�Z]�/����iM��*e"���Z��#6r����;�L���9��Xv7�j#���1���Q��ǺΕ������5�)[���h�j�i�+-�6��.��L�L;Л���������B�D�F Ho}2b<�s;-K�z
R��h"�zP"��/��q�&��c��:KYܼCI�_��7s�9���o>��l%i�-}ϼ 8���?Y��}ٹ���8TO��xÔ_��������CyW�f�tR�wX����K�Q�7Q�n��C���	�L�de���"�m���r°������R�wX��}�
�?�Xsp#HXD���b���#�a�x�Vx�%L��W��_�ړ8���/����,D�85Zt��= ��2��O�=�ͦ�I|{�0Lʡ;�¬pX��g��U-�e5��e6²��_�Ps+1���'���n`5�fK��0z�cUL�_��._0�+���LQ�.�v�L#�?�z�C���|�F7�_��^{ʓ��(%��A��7A��(�n��rs�i��<�M�AϦ6��.��L�=��gr(��������B�D�F ���*�;�Cg)�|q�4'���Xw�j�7���{�6�e���ӯIJ ��`y���_���e��� X��V�+�3q�bx�������t%>^�ߦ��|R%���(R\֎u�I��c��k��V���io����=�6��#ey��8�ib͠�Ԏl�Б���� �VL�(\LVWy�����Б���� �VL�(\^���>�Z]��.e���2J��`�љ����\���*��[t�gR� �ұ7���?�!���bJ���_��s�֙��)yX*�+�@��-��u�Y�KGAc<�p{�5�O�%E#P�u��� Sf��ƫg�T6����Q�u;��|B���r����ْ��4F��u�Y�KG�ξ������eiqb	��G��W+��W�y#׬��5�U��)���Y;e�iKI/B޾PscX{�X!,d=��¾ȼ!�`�(i3xjzӝ���I(͂��-����!�`�(i3��TBd��pS�*;q��=<�6>e��0�U+�qbp@�!�`�(i3�G�dE�h�����?uA|�d���{_8�Y��=�}�Vݨ��}Dq�f��mJ�0�6�!�`�(i3��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����;�jmT�#�,l����M?��y�!�`�(i3�2��}�������Ə��.A`��x ,��rQ�f�6l�}��}Dq�f�!�`�(i3mj�B��Vh�EtC�<�8
l]]y�1hPR����p�@�VҒm�!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f��Fr��jr��*�t"#S�K�.�w�R���y��q��R�E�i�m}66j�"Hs�w��0�[Je��0���*ܐb�m��v��z�Nc7/��.㟏��Z���2��}�������ƏCw�Hm���<��>��φ�?'�QW����GS�*;q܋�DKY��,Bp��S�HN��R��?�d���&������?fb��;_��8W�w��fD*�n�'��%Ǹ�!�U������,n/�g�.���ؑ悍!����م���R�{@�a��]��.e�����م���R7�j�2>����?XW�~a���@=�y�z�:k�_8%ӏ��Z���G��^���_--���g���R�?KYC'v�����p�*NiUL��˱�����?��řA{���r��H�+#N|^�V��	��yVoJ���'�{\�.�]}��=��YV�v�\�b͐�	}�@�w��˪?�-���ei�^�̷ؠJ��:����3���F��&tS�D�]v1�_ُ�����Ə?X���V4&�]Pn��J�:�_q�pWS�*;q��[�9w?�J�^ⴠfH {��u��]'\gWg��	�Z�kfc��2���80}}��*�H�RtV�^���{���#�0�zG�������&G���y��lDX�t�VC��b_X�XV�b�z'hۉ)��d�7�qĝ�\ NhtiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3���9���LQ�/8^3ZiY���Fz�΋O�»%���]c���HE4SG���Z�����T�R��!�`�(i3FwZNE�&tS�D�'���Xw�j�7���W�6?���_--���g|�m�ߕ�><���@��`.��53���w�@V[Z��.�~�5�Q�d
�:qEp}{e�z���sȸ�"rR-��ټs�  ����'Z鎬�������(����.��$��Rfł��kS�*;q�ց������b�Bϱ�mj�B��Vh�EtC�<��R@��"����Fz�HN��R��bP�63Z�t<�6�Q=7�A��\R��c���鿡�t����>3���w�@V-���,W������0�� 7�J�[|�m�ߕ��:5A��p0��l!���O�D mWN��\ Nh�;�P�t�50��l!���߸��S�ȌX�f�βB�.�g3Z�j5�{�S�g�E���dZ�,+$\�M��
,�B�UԊ&�!�����������@�L���SM�O��N� �P(����\�0S&",f�e��p�.������+Z}͐�	}�@�w��˪?�-e0��Tqmp�AJ�e�$��8y�Ɋ����Z��d�G}%��Ď��J��QCT�"�x9�¿Y�����Uغ���'3��	�.8��.��r
���иܖ�C�?�i}9]���Z��!�`�(i3��`!�r7��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!q��V���'�Pp̢���>�W��*(��3H��ieLb)�5�o�' ���@�0�0c��L>�W��*(��3H��ieL���]Cr$' ���@�$� %7䨉��%>�rG6j�"Hsʆ
q�8"�@��v{�G�U��k":�ct�0��3��O	�T/ k�|6�8�a"�/A$���Z��!�`�(i3��`!�r7��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!q��V���'�Pp̢���>�W��*(��3H��ieLb)�5�o�' ���@�0�0c��L>�W��*(��3H��ieL����A���_�3�|�.�>���@]��}Dq�f�����,�ǰE��C$�����B���'�綅������>vD���&l����$�<�F�q;��|B���r��������o�a�NO�*b*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+SƏw0��N�ijR2t�N�/�ڂ�nF���<�W�.�P�	��
�Q�}�.�g3ZQ�ͼ���ݑ4 ��3]�D��NL�G�
Rv��5*s6=��GZ>.�0'j�j�Jy?�d���&��ݚ�Н��9�|���l8�48�{.S�����g��+˘\5���jmY�wΦs� ��6��.��Lj�)6)-
FkH���8ч����B;�T�dN�<@Iv��nt=:��:5A��pw�R���y��0�J���Ė�b�����bx�8@�@�	Fφ��<�6�@a� ���N���������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�SƏw0���iD.l^S�ñ��̞�{_8�Y��=�}�Vݨ��9��H+�o~葸ֿ��OY'�E�g�������(ӈ���m�r����̢k���"��w6�0��ɗ��zi#Y)M���Fe���2+mxH�qV�"T���7X���c�}��
�t��T&���LQ�/81tSjv���'T���+~~!"s�(������6��:[+b��'�Pp�G^����Ă�\���tl&�� ���?R ���`!�r7q����1��,H/��HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�ȌBt�u[6K.�yў�о��#I��O0Y�6j�"Hs0vZ��ҹ0�(j��0���u���k�B^�(��E�1�����2������<�b���]F���2������<�b�5L�T!t���m l�o66����~�"���D��j#�{D�A�W+��W�7�:t�?S/��j�VD"�7�,��n6�o8:4�I���c�90B3v�A��8����z�:Fa�7��-Ukc��R2�e��b�uz۴k1��˲��y��lD=�1��*�
�I(͂��-����!�`�(i3�ٻY84����<	s/�=Â��'e��0�U+�qbp@�!�`�(i3Z��}	���C�ݥc&�̢����{_8�Y��=�}�Vݨ��}Dq�f��^{T~H���^a�nu4Bޗ��jw�	���ݚ�Н��po守�u�,l����M?��y�!�`�(i3;�E���� ��H3�յXg:�$N��GZ>.�0~�{ ���ݚ�Н����y��lDU�n�X��z��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!�`�(i3�iڈ(��֟�z��n� ���?R �����⪂!t-�u	D�&F�WAM�Q��\@
��:�)�<�����⪂!t-�u	D�&6���G1�Q��\@
����G3҇
!�`�(i3�I��Yqi��,�S��@/�uw)"/��=��K�R��K<_8 �B� �b��!�`�(i3�� л�U�~�vmȋ���OH��c���鿋�E~��k}����/C.�L:,�s L�Zl�W��{��]�L���/=9'�����mC.�L:,��i���A��ݚ�Н����y��lDU�n�X��zq����1S�Д_9[�l��a+Ĳ
�),��Tt�j� �"�m���r!|�α+!�`�(i3,�u�S�(+� �e���5*s6=��GZ>.�0'j�j�Jy1tSjv�!�`�(i3�B�.�4Ӭ�P8��PS~�Dn��i�Q׭n�L���/=9j���)��Q��\@
��:�)�<�����⪂!t-�u	D�&���A3�Q��\@
����G3҇
!�`�(i3�� л�U�~�vmȋ��OY'�E�g�������(ӈ���m�r����!�`�(i3��A✵0�ݚ�Н����y��lDU�n�X��z��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ��:5A��p!�`�(i3�iڈ(��֟�z��n� ���?R �K7͍��|��W&":�ݚ�Н��� л��5ߧE4��!�`�(i3��Qѳ$G��A0ok�®� л��5ߧE4��<�6�Q=�׹�%G��^���j�VD"q��_N���Qѳ$G�;��|B�6�'Z����Ct�g��^l�������A$�P������5d�`UNP�{y����:�*" �`�r$ɓǃl[�Ƶ�1tSjv�SƏw0����H:H;��=<�6>e��0�U+�qbp@�՝� s�#04~B3��������h��`�����y_�mS8<�n���F�P�7��S��h��d\�����l��=�O�-v�*_�mS8<�n�ݚ�Н�!q��V��hiLi?֑�3���iD.l^Sm4V2�@o~葸ֿ��OY'���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��'�v�|u�o�����V����d��U���q�z�#˭����A��/A��CQ���\���Z!>�-ᴘO��8e0��Tqmp�AJ�e�$ũ�R����yDƶ���W��d;.�Rɩb(�7/ h�� �)Q���k�#g�k���:��Ɂ�]�'߭`��@_��M���o��_�Rv�䩲$���dS@Ɵ�od�G}%��b�l)�=����"sS<�0�zG�������&G��'T���+Ho}2b<��8�.-Mb_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3���JQ����c�0�=�8�tw��~~!"s���̰'0���]ԍ6�!,�:�֑@�VҒm�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�\;/4ҟ��,���Ъ��}H	��*����,�ǰL�[��V��%am�m�C��߮˻��b����ق��`� a���{֐��<ͯ�G��R'),��`�a"��-K8Pv�f^�fǙ#Y\��?�l~�U���� G��n�r��<� �&���=�k����D���n�)�<ͯ�G��R'),��`�Սl�È6|?�d���&�#��`*�Z�u�x�c�lR��~�IX0F�MV�ҁGG�.Mm-;�C>��Ӛ<lȕx��H����Qw�c4~Nr_�mS8<�n�ݚ�Н����JQ����c�0�����AIe��0�U+�qbp@�՝� s�#04~B3��������h��`�����y_�mS8<�n���F�P�7��S��h��d\�����l��=�O�-v�*_�mS8<�n�ݚ�Н�!q��V���팣+��F��0vP�E�9�|���la��g�p��_'&�d�'fU����"��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�"v�(=�@� �-k��!�ˢ6j�"Hs��'���5W��.�y�Ts7U�] �Vl%���'�١�31C*e�r�_���w�BVn(��ҫ>��?B6o���J�$��F���A��S&ϊ�`�y���z,3���� k�U�y�3:`��7.C=�����9�� ���?�$�i6^�W��2��~w����[KX��q�}���D���m��g�k��"]J,�O,��MR���V�^9/�)ļ���ud�H�V�܄WD��|���l5R?}�b�k��԰�/"��nH�W�v�7�� I�����.��4�F1����jaս"���H�V��=�WK=Z�B�
���}h8oS뒐ȋ?4wK�G�5���7�E� �y]Xg��n�����wx0�<��w��Qo���H6�կ��\��D���&҂��j��-�����#�Y�Cφ��<�6�@a� ���N���������y��o��7�;�jmT�#bs��2[�a��o���H�RtV�^�#~.��,��tE�ӻ���+.S=dN�<@Iv��nt=:����q��{d�ƥ�졪��'DV���b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3���JQ���8�0�&a��;��]�!��	Ǹ�y85���`�8Ә�!,�:����Yմ�nJ�|m��g��U-�e���+s�Kv�ء�����6屍Z鎬�������(���0��B�YV{��>���|Ƅ{�6�eυ���K��k/��m#��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�"v�(=�@� �-k�L���|���A��S6�w�*u��S���m��+ٰ�Ř�h�f�~�?�M"`h��@t�iZ]XF�hx��G����Tkd�_Ji�];���Q��\@
�Q �H����]g,H��vє�&���X����?����O,87WA��s�E���g^{ʓ��(%��A��)�^�\�E	v��o�1Ʌ�Mi5�'�@b��Oa�@��I�Y�K%-H�V�;���)"������w6YmC,iguGظ0����t�%�Z?�MZ�ʛ�z���dЕ�ĦsW�0�c��,�#���@��^{ʓ����-�����<ͯ�G��R'),��`�K����F?�a�x���x����A�l$�+9@[�_zβrE��g�Hbc�m� ����\�Q��4b&��K���w�����z���o������,�ǰ�QCT�"��I�N	�7Q�n��;:��_)�:)f�����9x��p��;mQ�MM
��,=�GdC�b�>y�T�.�~�k��D����팣+��A�׭�%*be��0�U+�qbp@��-��~U��j����J�;����<�����;�)R2�bP�=�ƛ������CyW�f�t�}+N_q��(R\֎u��Vv/�y��{pxʟwf5��F�$N!U�t|�Vx�%L��W��_��MM
��,=�GdC�b�>y�T�.�~����`���ƼP��d�k��԰�/"��nH�W�q3��+����/���	0xǎ� 3�kM=/[�)�������sP�������tw��ĕ[뜗��,�ǰ�ƍ��i����E�p�2W���R0?�@�|��Z鎬�������(���R0�����%��Y���#�����.��4�F1���Gb	l�%T�#�S�� n`Ip�\{ف(�7���<��Y�&l������8y�Ɋ����Z���F%�X�ԼQ�}�p�?7P���`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��?KYC'v1��E:z�'�=;v�����Ə*J�X�$��c��GlhŦ�.�g3ZrZ�0m�\�S��u���F%�X��/����7Fk����PqZ�o���ia������v�h�g��U-�e a⣃_B7�}�!���u��g��L1��E:z�'�ĩk(�CQ�r��H�*J�X�$��b���9C�.�g3ZrZ�0m�\�H�z��.�g3ZE��g�Hb麭�H�κ;q�+����Mgw�� 
~�F�,���XF:6/������,���eFz��^�̷ؠJ��:�����0c/��kk��o������"O��_U)�<�&#R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G��^��jsrCm�k�:��=#��9f2Pih{Ø�Fɝ�\ NhV��	��y�� �P�qN�/9ݦ�R��X鷴QW�w��fD�W�_����Rr������%�<�$