��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����i�'������\�-ǋ 4�i� ������[���a�8%`��4�s�6�XAoeuxLZ�#8�d~O�GӔ�<4��ˌ�ň��h��=i�@x_\q�jB�Fg�Y씤`��p�܂aQ�"6�l�:���3��>�U���T���딣0&_���X0���2|	p��rw@	@us��Nิi'Y0ii^sZ��yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪ��v���4 #e�l(.��>��'��E����F+��T����g�"�xI+r�� 0�D�A�f�mX׌��1w�J}�tGvH���O?�
'���}@��r���7�H&�Y����W��ĭ������%�_�~C�8"��� _�<�4SJ�����������Jw�C/��!��}9���S岦�%I^��������裐d5���Xf/vA�VG��ΊՉ���9?�\�N�{}�=�v��}�����Fz�!�`�(i3!�`�(i3���D��ܒ���-=*�ћ�Z':����"� _�i��i���5���6*�t��L�kq�]!%����<�p��G0�=i��/$�ߺ��]ַOk��!!�`�(i3!�`�(i3*8�2�z�����b/?�8I.���^r�b(�c�ܲ��F�t�Z�f��I�P�Y5�����c�o+��L�/�~8����A�߲wb��� ��WM�P[����(,)�=!�`�(i3!�`�(i3�>L���L�ɚ5���x�[�%���%���=���pw�ۢ2��vR�J���}���	��!�`�(i3!�`�(i3}�E%|0�WJ�Slm�m��}����ܲ��FC�����էam�X0�(�'�I�i���^�w\_�Z_!1�2t��d��Z�����d�*���Fz�!�`�(i3!�`�(i3�7>�����D/͘B�5�35�#� "�q=i�/�J�0�)�u',�G!�`�(i3!�`�(i3eI �#��I_h�R$:7�����m�e6�B���k�c��`�	U����f�7U�i�#!����P�>+�va��2u<�F�x��_���RQ�
�0��,��X!�`�(i3!�`�(i3�f��mt�5̤뢲�
�7>�����ǚr��y�v_4~�X؟�r�u��Q��@YO��<$e|����w'��1�:�Ω�s8�R�	�}����i�'������\�-ǋ 4�i� ���������	x]��/$��x��~篟|�Q�M�u�cX8N_�=rџ�_�v%����E�)��|������\�4�sg�oXx��U������ՈĀO��w���9*<��*{�ۤ���*c���4�a6�N��?���\z-��EM���
+����rx�]�V��\#O���o�x��`�|>���P��f�>�٘\Ε���}�P�������pC-��h��☂/x+��s(a�L�"�,�9�{��2$6�sI�حЄSZ�h�5L��p
� �AH��1�����m'���h$��ޝ�~J�,.G[��	�F@�4%�}����b�+gobQ�el���V4zm�!=�y����h�}?�.�10�.�	�Z54�݁y�k�����}/��)
��4<�h=Է`nӸW�{|����u�	H�N~��v�kC���r�O��C��0��]�)හ��I��pg���P�A"KۙJY�7C��H���`\����~�/���3�+��RL�a)'r�Ӟh� ��I�;��mȨ"2c�P*�^�7C��Ho��B3�;T������v��㡝�r�O��C��0���t�J0v���I��3Qq�^U�|s.�!�zg�Z�$+�~c(�U���.�O'�W2�����`�f��ϵ���Ԃ�W�o�r�O��C��0��ד�̟a�,��I�U�߷� �9��0-*�&�!�zg�Z�$�H�`}�f���L�B�)�g��I��fP%�SyI�D���i����	x]�������7��Mv�9��a�{�0�!�C��jџ�_�v%�#���{��Hl��f�� ��C���)����Xz��BV�;,J�l�/���D��ܒ�L�}��B���s4y<le��^(hO�Ԏ�G�K���y�\�ʆ�In��t0�'�@ip@{,�����O�Ԏ�G�S]�����<u��w)�S��X3�������Φ�8ưc��!?���5"D7n=������{wÎeT�?�)h�52���,���+�k�8���҆�|n���:�o�E��Y�����rw�O�I� ��ѕ���Ϫ+2��z�W87"�o�9���1�r�O��C��0���df��/w���� �b��j3�w�>��SU��Pa�s��_;%v������J��\���a6�Ͳ
�3�K,��,Iw�)�D���i����	x]�G�Lm=�b�7��Mv�95�KP 4Z,�&�$�kyKџ�_�v%��"3<�Q����AyU��Z��G���Q��ȎC3	^Yt��m�ep����`�����F�*�h�҆�|n���u� �(�ⱃ�!�QD�:mF�'YJ�Й�m���K#Q��-�Q�\M������L���ڰ�]���]�����Uˏ

�2�ո�R@�2r�O��C��0��$�>��w�*��D����Ǳ����w�>��SX`X�B%�r���7ȓC�-`�e�g��!��x���� �"!B�������.�-���
E�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s���ħƿ�9c:��{~v_z�m%̼�{���_��w���C3�k�����ΈIn'�J�gs�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�ĲW��,)i/-�#�����ˉ�1�:�Ω�s8�R�	�}����i�'������\�l8������ea�;y� ����t��=l�)��%�0|]<w:����+�J�������V����(�}	g<��
��Knc���9?C�Ÿ�-��p��ڨF�:v��Q�^�y�����9��;C@����F���m¡B^`ٌ���i��؞�%Ah�%4
>��f���T,}��I�dp�S�5я�����0��zO�) ���3�ҺMC�^�.�]V����(��wl��h�,|ފ������o����[7�d|���f���T,}��I�d�p�[�d�G�@�Yk�.�
����>2�}���!T �����c�Y!�`�(i3!�`�(i3!�`�(i3!�`�(i3�S�����Z��L�*P{���2����$Y��C�5����*E�eNzL�lS��V0Ӹ��QC)t88���wH6�x�{�Z��{��R�wtJi���M�C2����m!j��Ę����@~��,���@ݎ�T��ߞ�����i����D	��U�q��w\F�]I�Dd2�Ĺ�������w��Ń�S�16P! ��:v~E�)d,w0��tb5��Rb��Y�W��u�Y��2!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�*�2߄�ѹ��p};�B�v�U�������T`���Ot�rZ�?ђ��P^(�ՅG��u
皲��+�J�������V����(i:o����|�������)	�8V���C~��m���4X%���'�4ɀ�i�X!�!D��(J�f�'��q�S<MC�^�.�]V����(?��I��I/N���{��c����ma���q��w\F����_�.���r'��˝Sz��E�4.@���u*K6HY_���P[�z q�"MI<��fҾ��9�����?�!�`�(i3c��Et��q���U�ЂDa��(���o�d�c��Et��q���U�C#/<���q�VP��@�����ɧ�J�8�J��	��	Mk�r��|g�Y�'���Xw�#�K)���J�I���|g�Y�'���Xw�j�7����w�K��ݑ�][HW��W���֨g��U-�ee�@Rv����my$�N��o�/���;vwdI���<�_�r�)�s�ި��o�t�����sRt���j��\w��0]�o�t���Pm���7G#+��\w��0]�o�t����L�u����j��\w��0]�o�t��3�i����j��\w��0]�o�t���ԟ'�D���j���0z�cULy`�_I�v��4���OTWRdr�Jbk-����'�\�n�wa��>���g��U-�eaԗ5��C�����/��]o��in�m��+�<4��ˌ�ň��h��]�F��������Ah$��>2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc@�����>P�2-i_\_��� �yz��$6�D��L���_�L����\�Q�u|v5�*�.�z,yZ?�X���!�G�Ḁ��Ʌ�Ě&/�7��6o.|�^��
�>IÙ=�Hs�$�[�k-�E ����n��X)r��!�`�(i3x�]�V���Ù^���Ah���l�-��;���,DtL�㎭J,�t`N��B�:��c���'���Xw*���������@-=�8��"�7ϖ�|�������;�71?9Pjp������PN��a(􆿳��ȡp��'���Xw�j�7���7>�����ǚr��y�_��wBW��8���/����,DU�m#j[-d)��5(�套�qD0�f��p&d�@����gG{�bW)Yq����Cs7s�9���o>��l%i�-5�e`��9֯���,��1�k9�Z鎬������_�,���R�A0^L S������Q]� _�rs�i���`�M�	=̞��>�B^`ٌ��x�[5��Z�8���/�,��Px��H�u$2�Q����4|����߳�wM:�rQRт���+�J���q���U��@����gG.��U3�
g�YӅ:�7s�9���o>��l%i�-�u��Y'GZtgQ�9OZ
�@R	~��Z鎬�������(���/��A����Q[R�7�
�CӞD�߿�wW����8�S_&Z鎬������_�,�e)����|
T�W����Q]� _ό���.�}�
�?���U�R^p���P#�d�٣���N N�S�dg�W�p᢯��0�F�?�'���Xw���,D.5�����O���Wśy��n`5�fK�\w��0]b!��u�ì�u"4�"�,�>E����\�v�g�W�I吱 �']g�׺�&\VI`,�ϖ���~vJ;��	�yE�Ss�x-��A%X�z²���ʓ�*Aj�I�e���_�$��*�yW��Xi9�
�іm��U'�k���W�f����ހ�Fhʢ!�5��=l�U�-��#x�۾����!d�h��<�qƂ�$�������i��O��$��Xo��ߌ;޴@�,ԯ���gn"G�q�������b�3!^�3�@ym�-f:2�	�^����Ћ�l�Tq��W-q�C<{�uig����V�dN�<@Iv�O�ȕi�l=I��nȑl�5��̄qbqlФ�vt�q��gbb˸xZ鎬�������(����\\�*�}!�X�V0Up�rP��O%�ud]�M��+x�r����l�©�]t��):�Z鎬�������(����N=�[��e���ZF��ֱ�q������m�q��|�1��TZ@�6��7�){`4�2N��n�`�*�������r���Y�{'%s�6F���y�b.�hFd=��¾ȼ�u{*�C<�3�@ym���Ζ��1tSjv��37y���� ���30��w�w:�;�jmT�#,��T�����\_���/]�l�����&G�q�9�ͭe���PO�my$�N�����'�ډRa])n#���r������vf�<�R�{_8�Y���0�-��Q����ƾ�x�\oqv !�`�(i3yY2�̾���U�;��tS�$bnNfĉ>99��A0ok��[p�#�_ wgf*��$�Q�����S8�&u�η��.�[�X��=�gw�⽒���n�����:=�e�)�ή@���P��� �Uj�.�B��0�9�@�`���}Dq�f�Goj ��6^�h����!�`�(i3pı��0����%�m1%�Z��3��w��\�W�ƍ2���lĵݓ�W����l3]�T4�0 L?ஹ�%�ԟ����U��ݚ�Н�(*�O�q�ͯ�*�d�[}�N�`2���K����A0��s!�`�(i3�u�24��&~e�e��E{��h5���՜����|e"ʁ���MյX쯢86�	Ղ�I8�y\��S��z���wb��Z2!�`�(i3U /숇�]�	bC��<-�;S5b	��T�.�w؀�CF��6��� m�#;[��U젩`#FW8�	����C��s;��}Dq�f�G�&ց�*�=��
��P�n���}���S.�3��"Uʡne�!�`�(i3pı��0��Y�]�q��c�Z��3��w��\�W��@�����ݓ�W���D��!~�4�0 L?ஹ�%���EXc=Sq�ݚ�Н�(*�O�qm͈���߀[}�N�`2���K��m���
`��!�`�(i34r2p�jg�&~e�e��E{��h��^9�Ƣ���|e"ʁ���Mյ)n�B�D�	Ղ�I8�y\��S��z������'�!�`�(i3U /숇������<-�;S5b	��T�.m�P��/A��6���r��(d��U젩`#FW8�	��2g���ܐ��}Dq�f�G�&ց�*�la�T�H�n���}���S.�3��7�E!�[!�`�(i3 |������if��Y��Z��3��w��\�W�ed�N�-�ݓ�W���	�N�M���q�嘝��ஹ�%��2V[���X��ݚ�Н�AL(�z������0`�?�JY�)�q��ڍ�����a�"��6���@�HN��R���ء�I��$�S�in�Ye�ήT�C�5y��;��d
z����YUr�(��z�j�Рe����:
1���Ʊ%5�����꠼*d�m|ag��6����?�g�˖���R'cf��i�X!�!D��(J�f�w]�IB[�)����]�5�O�%E#Pw�����A�#���Q�XS�Д_9�	5XYUʛP{��Lג�Q^�MY:�6���;b��g��U-�e��:���j�D24N<I8����\.W��/z*x�n;��|B`q�a�i��E2�DZ��(Ɲ?��$;�Ղ��5�ʑ�(4K�I� ���F�Ҡ��q��É~�nJb�G �!�`�(i3�3FV�J�3�gI�f):������$��z���q��l.�2N��n�ܖ �&��ǳ<��C�
�rA���oq��WX ��b�FP&;Ε^���N>I��WJ�jݭ�F���%,�������;���EWrAԢ�a\蟧��T�j�c��\�v���+x�r�\�,�
Y�>傀��E����F����o<rS�b�8Z���oگ��r���%��Q^�MY:��H<㕕ѿK��#�$����v���$�Qu�N�#f���C9*�¢�L���`H�j�7���7>�����ǚr��y��CyW�f�tR�wX�է2N��n�S�/��8'�-Q?9������5	�3C���_�����8-|�D��Xmt�=���3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l��@;Z����q���f�e�x��w����֯���,mk��L��x{^4��*m!�`�(i37�%M���6Y ��؟�r����ڵ�a(􆿳�Εq�8!�`�(i3�Zj���
�7>�����ǚr��y�%�!��U]�ߍ�2d��3џ1�F�Z	��;���P*��g��It\$�ݛ5�CN;���P*e�{�W!�`�(i3.$����0�*��D�x�=l�U�-kO��u�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'��a�}o8g���?�!�`�(i3�k��^�1Jbk-����'�\�n1���R��뷅Kn�;F�Q��s,�~TM�e�w�G�;��]�I�h��\�
oOݎ�T����U�s&����\W��N�!�`�(i3�Dd�\���؞�W�}�:�c? ��@2A^N�]|-&vY��;�!�`�(i3���F1������$�ӿ�F{ј�^�ݚ�Н��Ra])n#����m?�V?��?s���9qj�xm�N�e�{�W!�`�(i3"(<K�'PyQ���4��}�@���_rS�b�8Z��W�6?��O�M:R	�گ�����ݚ�Н���6������S>�D]h����yQ���4�uE9�+��!�`�(i3����١�$�ݛ5�CNTף�[t�����������G�R�u��r��!�`�(i3��>��lJ)�W�=�k�Ҟ�#�>�L��n��p��b�Bϱ�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'���Q��\{9
Cj�R[z�!�`_q�!�`�(i3$f��_Ub�F�S�1 �����l��#�X��C����Խ�TЃ�si�ݚ�Н���6��b�8W�wo_V��U'��Cq_c�!
�T�r�5�!�`�(i3��jVѭ@!�`�(i3�Jo���jQ�kŕ��QzM#��m�<�6�Q=*qm�U��g_WԽm`�P^��ݭ%�?�p}iBy��R<�pc!�`�(i3���F1������$�ӑ���n,��>]��e��^���!�`�(i3HN��R��bP�63Z�t!�`�(i3�5ߧE4��!�`�(i3�u��A�0�Ή*��a��2S����Rq� dr�+6V��\"��C�/�y|2I��jsi��3�a/� h�ҩ���6��b�8W�wo_V��U'��Cq_c�!
�T�r�5�
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�g��ޏ�Jw�)��b��6~����7���ċ�Pm����5�:�ဧ2N��n��|�'豪r+f��"�r�Sy�n�yLjn�=m�"�2N��n�[�hŽ>��3�A���u��s$y�`�U+�PAN}�m��{�`{��U	]��n�fyP�?��{	1�Z8[iI9�o«IX0F�M���&fy,�3 l� ���Aؠe
�M����'����u��r��]�.�,���9z���@�oS��ܠ�a�,��
�T�r�5��po守�u�tu��#Ǽ{ڼ�`a3DGi�s^z�5�H45���֔;�K�Ѿɪ�K<�����?�~��|#HK���\�A'YE��"� _̸ ���]�0��Olz!ב}�bg �}�7��H��"� _�W�}A]�)�� h�ҩ��o�t��z�
1���;n��뾦�՝� s�#���k$ �o�t��z�
1���;%��v��!�`�(i3��J��Gv�;���-����!�`�(i3�R'cf��i�~�B՚��Ʌ�Ě&/�7��6o.�@�2�2r�ݚ�Н��{�6�C������n/��dc�@c�����h��}Dq�f�HN��R��Gu�"�0����%>�rGO�D mWNHN��R��bP�63Z�tU�Q��$�n�'�Jh$��Ȝx�����\�J��w�w:�<�6�Q=�5//���"� _�W�}A]�)�� h�ҩ�V6Y��@��֯���,��e_c�?D�8��v�0!�T�ݚ�Н��o�t��z�
1���;n��뾦�<�6�Q=45���\}9t�td���5U�Q��$�n�'�Jh$��Ȝx�����\�J$f��_Ub���uQL+��φ��<�6�n%���H�|���[�: ��뮭tn S�������t�T��?E-h���U���e��_	�Ƽ��S�J\7fF��v��T�#��[J�;��ܿ����qD��=a�^7�1tSjv��m��
��m�a�gPM��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l��3Ҝ}�u[$�w)��
=b~*��s��0M�Ŷ�Eʨ�`N/��R��3����'��a��o���H�RtV�^�9lD��XH S����<z7n-��86�aI�[��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�����RCT�I�N�A$�:��EVu2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϓ���T�����^Lļm����7���eo~��.}�՜�����GU��L�z����:2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcW
��0�X���:3p�k����F��o��_�Rz���n H ��b�FP&��N�T?w�W�E<HӍ*"v%)��2�����B^`ٌ���+A�J�ʥ�n2`q:Fa�7��mךBo�NX���:3p���IM��P,���^a�nu4Bޗ��jw�	��9gp���mV�I>1͊���3-��g�MSG~1tSjv�U����ޚ�W�o]��e���Γ8�dKa�����Q؃�L��r|����$J�-��^�����H�����?�@,��V��J����(�ߜ1�fR��}���;�P�t�5����$�����F�z�8#���1A�QzM#��m����y��lD5��ˬ�d`&c�'N�jτq"�;�A�b��Q���N�T?w����L1��3��`��Mupͪe�>Ht�u�Ud��:Etj�/��@����	X%+�=�x�N�M��*�8��S�҇�8�\��(�A�Q*�I+Z����]�w9"x����l���^�֪P�ꜯ}Dq�f�1��3��`��Mupͪe
T�W��d��:Etj�/��@����	X%+�=�x�N�M��*�8��S�҇�8�\��(�A�Q*݇\��"4���]�w9"x����l���^�֪P�ꜯ}Dq�f�1��3��`�����
��A�IS��03�� <I[��hg׸�� �?Ct���g[��p����y��j�ɋz�����#~胁T���AZ���ϛ?
�ǈ�MQ����ry�茴�������������F��帵dE�[dB~�S;����Z<��A!&�2����M���CO|e��߬�x#=���c���9���G��_�t�^��+�"#��̒aF��&�z. �G�4f�e"ٝHN��R��bP�63Z�t���F��O�\E�W��4bmךBo�NX���:3p��G�tM쇱|�G��?��Ϙ�q����#����6E���ΐ����GW���6�o8:4�I���c�90Mj�dL�{y����i�q,?5qj�����)�_3��Q�dxjzӝ���w3��׍�&�U��f�tl�:�K���(L�^5%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�`�zmj�������XRߖ��4!��1�b$`��g�d�H�RtV�^p>��C=U����]��"��ӌ�r���%>�rGO�D mWN;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���!*��*8M*QfY�"Z_�mS8<�n�ݚ�Н�4F�M7�ũ��&�X|�/��kOTfĉ>99��A0ok��HN��R��bP�63Z�t�5ߧE4��Fr��j2�d�6?�;D�Vh�����"��3y�ܐ��H�ǒ��~Bۧ��߿�wW���Z<��A!��jVѭ@!�`�(i3�2 /��u��������[`&c�'N�jLm�<o�̍�T�t!�`�(i3!�`�(i3՝� s�#���k$ !�`�(i3�4��������Жm�᢯��0�Lm�<o��G�#����᢯��0��ڎC�?ΔA
i�eL!�`�(i3!�`�(i3n�)�� �g|����x�~c��0���IX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>�j�y��j}@?��W���qD��=a�^7�1tSjv�� �@[�鋽C�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-����;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���!*��*8M*QfY�"Z_�mS8<�n�ݚ�Н�� �@[������4Yz����|e"$f��_Ub�F�S�1 � ���Aؠe
�M����d��-��!g��J�s��z�
1���;#o�]�ʄ�k�q@g����Z<��A!��-����!�`�(i3"��
%��v��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M�+Y�6R��j�'l��@g� BO����U��)���Y;e�iK-pm!9�>��n4s1�U��B��-��8�2W6��v�����r$ɓǉ�.y�U=������&G�l�de�����$�a���NM���*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3����,����0�|섃Va�ir[��l�,t���H[W?x��w����]�Լ�c�G��Hb� h�ҩ��l�de�����$�a���NM���fĉ>99��A0ok���H�����<Df��Eʨ�`N/��R��3���:
1���Ư����z���!*��*8M*QfY�"Zg�d�H�RtV�^J>zߋ��>[;\v�a��ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}���$�uG,�د$�Dj9�J?�����A"�S	��1�3�����+�}�`��:Ŷĺ��}x4�Pe�I\��Y�tM��楱�o��_�Rv�䩲$����E)e|A��`���φ��<�6�`&c�'N�j��v�����r$ɓǉ�.y�U=������&G��(���0���;	ȕ?�q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r����#�a�Ą�ԬQ����5��t�	���QC�ڎC�?���> +�S�;��ԗ��8k��.ͥ�H�RtV�^��Ϟ4�>Ht�u�Un��뾦�!�`�(i3�5ߧE4��!�`�(i3?��LST�ed9��a��o���H�RtV�^��Ϟ4�>Ht�u�U%��v��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�Ms�Uo����N6-	��6<���{k�˖�x�󢯖^��'�ZT�����sz`F���.��n��܆���M�,!hޖ�A$�P��O�@י��2(��T�gu�#��nt��F�z�8#�b9���:&�>��s��n4s1�U��B��-���忔8l{�]&"(ShT������qD��=a�^7�1tSjv�œ&|�9�n�o&uL�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^.%ĩ.u:�J��I�s�(�ߜ1���iB��H�RtV�^�0�9&،��F�z�8#Ҟ�#�>�L��n��p��b�Bϱ��>1J���ƈ5$YaV!�`�(i3��jVѭ@!�`�(i3�����i��J����[���G�����Gܘ���a!�`�(i3���F��O��ݚ�Н���#�a�Ą�ԬQ����5��t�	���QC�꠼*d�m�d��-��!��b�38ܽ)f�X3G��'��b~*��s���v[2�����xQ�OO�뗛QLm�<o��w��+-��,�J��f~T"�lġ��j��h�j��ݚ�Н�œ&|�9�n�o&uL�״$(�>g�
�:qEp�;�P�t�5����l���a��Bަ.ȇ��_�mS8<�n�ݚ�Н�œ&|�9�n�o&uL�)P<�ܓ�Y
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�z��O�������������m>�G�\�Y�&[R�V&H� FMsO�~�fB��t|ql�osZp�W���
�$������%H��|���2,bK���ŃN�����U��)���Y;e�iK-pm!9�>ֱ�q�����ѧv;�?�@,��VJHn��z��r9�3d�G}%����3f���L�yE�:�.�N�������a��r$ɓǉ�.y�U=������&G��೹�C�A�IS��[;\v�a��ƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l�鑴HH��"�̙	,N��>�s�,�H��-����!�`�(i3}���yb���}�@���_rS�b�8Z�AԢ�a\�2}$#h6������t�_��ݚ�Н���jVѭ@!�`�(i3}���yb��-H��.�����o�����[��l_HN��R��bP�63Z�t�Zj���
���+1�;�.��1��!*��*8��!�qgy�`��vN	���QCLm�<o���(4G��>��L���?�@,��V��Q-s�H�RtV�^w-)Sz�M�:�.�N������4Yz����|e"$f��_Ub�F�S�1 ���p`-�F/᢯��0�Lm�<o��M?��y�!�`�(i3Y��8>h�|�Ȝ���q9+t�}�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���U�Rdd@��2ʬ;}it���U�R��>qO��\��Q1�dfC0o�4��F�悠A�,�v�E²�i��z��V�6K�FX�pΌ4-��FB~�S;��ZN����6�o8:4�I���c�90Mj�dL�N}�m��{|�v�����G4aL��zL͊�q��D2<�4j��`���φ��<�6���U�Rdd@��2�2G�,��R(�U���e��d9=���u��r��Y��8>h����z��q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r��{���v0yfb�YL��&\VI`,�i-W����� h�ҩ�Z��JP���K���&��N��Ưb75���J>n�	G0��p-����`C��O9�՝� s�#���k$ Z��JP���K���&�9�ڟ,AX3�T�#_�B�ݚ�Н����F��O��ݚ�Н��K�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir=5.B�����d��-��!��:28P����p��ݚ�Н�ըa��9�_�o�@^��*�f;��}Dq�f���Ě�����}Dq�f��#	�Bj�A�IS��,ܓh�,������&G!�`�(i3��U�R�ܬ�mо%��v��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M�Uʮ�V(Y�$��fG�aН$J�MF��(�[�o��_�Rv�䩲$����#��i��~�26��\;��B�lXm��G��*IÙ=�HV%~YqsوiI9�o«IX0F�M�sݸ�/�gxjzӝ���w3��׍�&�U��f��"�чE4�]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�.%ĩ.u:�J��I�s�(�ߜ1���iB��H�RtV�^U����ޚ�W�o]��e���Γ8�dKa�����Q؃�L��r|����$J�-��^�Ra])n#���r����U����ޚ�W�o]��e�����<+yj��x!�`�(i3�5ߧE4��!�`�(i3����,����0�|섃Va�ir[��l�,t���H[W?M?��y�!�`�(i3�iߎ���G�>Lo;c>��X�?��-����!�`�(i3u�st����'�PD�՝� s�#���k$ �B�'��a��;��%���b��~$�!�`�(i3���F��O��ݚ�Н�F< �ذVb���(L�^5#o�]�ʄ�ݟ�e.ama�`m��-����!�`�(i3u�st����'�PD����%>�rGO�D mWN���%>�rGO�D mWN�mJ�0�6�fĉ>99��A0ok�����F��O�\E�W��4b׏����Ӡף<�W�_2��VU(��z�j�:�h�²�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ſl �