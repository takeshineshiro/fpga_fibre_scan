��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�4��s�A�|Ԣ��g��B���������'QԵ���
yL��?� �~�ǴW{< &{�!�y�W�BE[��l+ �����)��(�@rD������tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�YZY0@ìO�tw:g+��T��٤�2[51g.� -��E�I�?g�f�$��P�`
5��*�z��Yk"1/���%	v3�.�z,yC�v�V�&1�.�<86�8m��+�����3�Χ��nEA����n���bN�<�B>p\�?;�+C-\:HBm��+e�(���n�JŬ+��M"`h��@{jϾn]��Yk"1/]���!E���VG%����@�/��(����5���&<˴m�mPۑ��X�b����@��q�©�lj�Ld눐�PF`H,�<��t��<vkS��1�:�Ω�=A���>�LZ*IV���^���������@�/��(����5���I�zI.�R7�$��p�S$�&�.�z,y�n|��ea�8���`8��xS�^���������@�/��(����5�?�J�Ń��ɖ�2i�螘c&H��Xj�Tm��+Ȑ E�������?9���Z=%�t��<vkS��1�:�Ω�>���U�_�4�0S�����x�M"`h��@{jϾn]��Yk"1/s�\"���a���ܻ�YD��bG�I�?g�f��Qө}�_g�?�H���w�1���i8�䟿��Px?w�O'�lR(���«�������d��M"`h��@{jϾn]��Yk"1/��n5R�%�.��.f\y㔪�_H��Xj�Tm��+�ڔ�wV��?��N��j�M"`h��@{jϾn]��Yk"1/+���鷦:`�'ࢯq@9kOg����:9�+�m��+e�(���n�JŬ+��f��WjCt�z&��ÃlO ܅d��2��̪U��֜��3�Q�^�y�zL͊�q��Y�tu�0�p�ϵ�DEG�p�P�� nU�IÙ=�HF���m¡���r��1�Z���=���u*K6HT�����Nb�?49��x#2���p5�}�]���x�]�V���KD:�}����L?V{��\G�Y����-�,�_��(֥�e.��xu	�>��l%i�-�M�g����c��Et��q���U�&��GE<�N�By3��<�]�!����M[��Ǣʘۥ<3���қ��]�!����M[��ǢQ�P��
S��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+�����
L'���Xw�j�7�����r��1�Z���=�"j���b7xY�J��ev�mS��0�
���)�*Y x�S��q�©����y,�m��M�5���.�V�k�J� VU+I��vMb��s��Yk"1/]���!E���VG%�[ b�����,\ަ�It�k\,آ()���;��G���9��'n�^0o_
-��[�����Kp&�@���k��l0��F��jT�����Nb�?49�����_�\G��4�	B45k�c��`��'n�^0o�!���!��x�	�2��g�P�e�9�:�]�^��'n�^0oM�D�;��-+0�l�R<�q��f�}��Gظ0���������5	���]���>����C�h�'f R�����5	���]���>����Cοƿ�d��������5	���]���>����C�?KYC'v�������|g�Y�'���Xw s4S�'�i��`�z&"hkIH*���>RTت�I7��-5��6��	���`y����ꢤ�Og�[N�&ѐ��(�
t��Y�{'%s���'���ը��_�\G��4�	B45��lC��U�T�\ ��Tǯ�!���#;r�����S��I�?g�f �H�Z����dn��A�.�z,yq��"�$"�N�p��G_�(����5���&<˴m�mPۑ��X�]�Xy8��;6aJVlO/8֩]=$���4�+|'�kP�?qNzL͊�q��UG�s���w¹��<d���<
DN��b9���j}8o{:�d�}Bȱ��U�p�[��i��i�����8�TPF�� g���t�&_���9��E����F�'n�^0o��ҕƦn+0�l�R<�q��f�}��?��[�<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����(��eظ��7�
BcyMu򔲊'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5��6��	���`y����ꢤ�Og�?�#B,�Ң�{l�f|�m�jp=�>��o�
�v�ξ����LUG���>��Oޏ��F˯�+)�"j���b7|#9���{k�h�++k&v�Iz7G#+�ǚ'b�t	�U���C��O]r�<Uee�,��3�L���&Ã�M�R�^Ƒ�Өg��U-�eaԗ5��C�W�T ��x���� �+��T�����h�6ؖ� onc�.�V�k�J� VU+I��vMb��s��Yk"1/�<4��ˌ��|��v���k.!�l�	�/�No`g	�ts�q�)3[�u8�����$G�yد�9�����~�����wl��h�)H��!n�'�\�J׽Z�ݽ;.p�7:SW�<�6�Q=Ի�弳$�.����~���kR$�kn���5���k�����L9��DUR�ߟ�;�Æ�MYi=�/M��%�p@Y�4Eb��ޒ`��`$���g>넽� �\Yy��M��(�K����!�ʭwV~���Vr�{r�����-N�'E�HG�vz��RxX��TԘ�H <8�k[p�M����G��u�c��Q��ݭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3j���T������q��
�e�~w�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�>.��̡��@��܊_�1���r�.v���t��W2�7�t`\���~��;�,!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�&�7m�3�i�V��wvf��q�d� s�\{]���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�z�-�v�k[�~�Z1~�g]�c�u��QF�s�����?!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD��� �oݗ����[2$L�e�(��0���N���z[�M�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD� ��*2�fNY��'�T��@�ш�ň6���D)9W �v:ι�Y7���&�_k�c��`�)\��FCR��]��e܅����
@{���e����q����؍��R��{QgkS�(!�`�(i3��%<�d�6�.�)��:�����y��j��k�s5=Ύ�9�j���B���7�F�ĭW�.�%6�<]"�:sNcbp��'�����U��ݚ�Н�`���*1R����
wL<65���Yl���#Kv���:1�#����az�~��c�&ck��K6�L+�.8%�����dN�<@Iv���a_|����ݚ�Н�H/�I��(B&�2�>��}YY�{'%s�&�
�0�pD��ZOU�g��U-�ee�@Rv����my$�N��o�/���;��6���m�XQ���z�+ N���>S̮�K�+EC�hHc�Ì49�����x�����s��l|�*"k���(ӈ��z&��)Q��!�`�(i3-Gb��F��E����Fv�Z��P,N�:2QYeƈ)P<�ܓ�Y���aR�!�`�(i3⤵�6�)�T<9 =��9�j���B�<Vo�eo���9�r7�K6�L+�.8%�����dN�<@Iv���a_|����ݚ�Н�ʅ|7@J=�P�:SôHaKv���ft�s� uƍ2���l�`���*1�I���`�����-VL�1���o�l����4�n���xǊj�ë��&�E���Kt�������qϛ�M~�ˇ�h��]�Hlu�����}Dq�f��H	EJF�dʀ�����
t��f"�	-7��8�r�%�
���lC��U7�C��zC@�D+���4Yq(����(p���	��
�Q�}A�����2�[<�!�� �w�;>cbp��'�����C��ݚ�Н��:#�R_��+�
�c�~��G1��[���J���T���b+}y[���S�fp�*x�$�Z�YBQ.K��]�!���\B��V���|e"h�wֈ�WI��}f����y���29��:|[%.�m�QA�Q* !�`�(i3H���L@�B�/�@TP3C6�HaDl����/	e�Ҏ�R]����pz�b'��nܰ��ْ5
�8��1�:�Ω�q��� �����_N���m3��> F����ȻD�ou�*Y x�S��q�©��'w��
�f��]�/V��X�f��WjCt�z&��ÃlO ܅d^�R@Κ�2���ei"�,�>E����\�vňu�,�s�^�R@Κ�2�l~�Uf���}��\�v�T?�7G|`�UxHj,��|��	�"�,�>E����\�vňu�,�s���2��̪U��֜��3"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3JHn��z�_c)���8���bg�1�Z���=�������b9����,����d���z���ߘ�)�I��<
DN�l0��F��j�q	k���A���������]c���H������i�=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3���D	��U�l>o��|�,+$\�M��wF4��0[����	��N�Ae�#����ꀍ!�`�(i3c��Et��q���U����?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-�|�)՜�4!�`�(i3v�ј�"��Z鎬����(��eظ�_--���g&e�l�����-��%Mm�jp=�>��o�
�v�ξ������ei]��fM?R�^Ƒ����"X��[��Q[R�7W����GS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l����G<�e��
T�v��1���6��	���`y����ꢤ�OgZ)[���F�����E��@IE�U��n�-�6��
�jW��D���M���R'),��`��{|*�"��i�_:���5�%]���a(􆿳�ؖ��d�I�� �:&�� VU+I��vMb��s��Yk"1/р�{:��'��F�N~Y�.�V�k�J��m�+��
J��@��ea�8���	�~�����F��mF�!؂�����%�}< V��,��B	hI�ˋ���p�ϵ�DE�U����E����F�'n�^0o�!���!��^�R@Κ�2e0��Tqmp�AJ�e�$�� nU�IÙ=�H��[[��Vp~z�r,����� ���3�ҺIÙ=�H�M�U�ct�:��RE��]n�� ���3�ҺIÙ=�H<z,Ҽ&�כ��p܏�<
DN��Q�^�y�zL͊�q���Vǃ����B�6�N@���k���E����F�'n�^0o4M,�����t������ݪ�򈟆�������\�vņ	N�1�.�]V�H7'�5�}�]���!�`�(i3x�]�V���	�?�ki%�7%1�e)s 3�:��)�[���6"�,�>E��4];ˍH�,t����t�r�hr�W�T}u��Q��L(\Ӧ�$�̎�)NC�lԇ�-{��E����F��j��\w��0]Y��
�iC!�`�(i3N�By3��<�]�!����M[��Ǣ�չ�Ad�!�`�(i3c��Et��q���U��ꢤ�Og>ݣK�6<o^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'��$Ι��o;�¬pX��g��U-�e�,���6+�mj�B��V%@��4��c��Et�Y�{'%s�[�&B�踫g(�r� k�|6�8o�`�_f>&�&i�"j���b7������[3���1�����}0xZ��T��B4׹C;�ދ���^�� �hi4J�jsrCm�k{��Kh��TD���rs�i�eB��P�ߘ�)�I��lC��U�T�\ �������	�/�^���E����F7G#+�ǚ'b�t	�U���C��O]r�<Uee��H�ʱˡ>mq7s̱!VkLs��dJR�^Ƒ����"X��[�'i�! ]���f�e�0
A���J��@��ea�8���	�~�����F��mF�!؂���������R$b��m�+��
J��@��ea�8���`8��xS�^������[ b�����,\ަ�It�k\,آ(&l������ nU�IÙ=�HF���m¡p~z�r,i��i���'n�^0o<H�-��*����Kp&�@���k��JHn��z�_c)���8�+�p}>&�&i�A ��E+���XP��Ȩ�wl��h�d�uY�ة�ʐx�?�'n�^0o4M,������2��̪
)\Y��7�ܥ��2��
[���p? E%n�/���i� � �	{����0�&�ͭ!�`�(i3N�By3��<�]�!����M[��Ǣk/�z�xEQ!�`�(i3c��Et��q���U�&��GE<�!�`�(i3Y%T��BPe.��xu	�>��l%i�-��TBd��pS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l������\�*P�I7��-5��6��	���`y���db�\EX@�/�M^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'"�C�ף�;�¬pX��g��U-�e�,���6+�+�uB;y�L�6yd(��(�
t��Y�{'%s�[�&B�踫g(�r� k�|6�8j��RO�I�1�Z���=�"j���b7xY�J��ev�mS��0�
���)�*Y x�S��q�©��ല���?�;��XCތ�; %���S��I�?g�f��r�F�5��I^ξ��ݴg��S�ZC%�}< V��,��B	hI�ˋ���p�ϵ�DE�U���JHn��z���z�O҈S��Ǵ��BR�^Ƒ��,ԯ���gn����fԱ@��2�F�P�F[`3*�!�`�����"IÙ=�H*.�PS���ct�:��RE��ʐx�?�Z�>)��p40�zɈ�UxHj,��|��	��b9����pP�o����y��lD�\r�q�{�؛G'���sR���<����ʊv.s/�B{�o
��P�1ߒg�A�/����<.+6J!�t���\�W+�[Z��x�]�V��;���Ӧ��Gjh�rO-�8j��zJ�	�;.9�(�4];ˍH��o��8�Ѵ汪#sЛ+0�l�R<�q��f�}��K�\7}�W,+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�H0l]��
(�5�%]���a(􆿳����^��+��%�k<�k��T<B7G#+�ǚ'b�t	�U���C��O]r�<Uee�,�Aٺ�Hᴕ��U��5�%]���a(􆿳�ټ*w2�56�M�g������{l�f|�ό���.���|��p��h�d �'���Xw�E�i�m}6*�3���f�]�!���D��L#�W�T ��x���� �+��T����5yi���FnBƕH�N�4�T F����ȻD�ou�*Y x�S��q�©���$Z�5�8z�E�^^������[ b�����,\ަ�It�k\,آ(&l�����W����\�v�T?�7G|`h�' L� U��֜��3�LH$��^��{�OF8%v@����fct�:��RE��ʐx�?ێ
7�\Z9�	��%т��!o.sG[�� �tS���}�#�ڊ<?@��[	J��;ι��QG�����U��7�ܥ��2�\Z�ؿH�j�\|Z��0[����	��N�Ae�#�̲�2�!������5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�^�9.�JQ�����5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�eן�-�Q�Z�pMݦ�l��-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0Tu�q�.:�TD��m�jp=�#{��p�{&l����_::���4�ˈ<�I7��-5��6��	���`y������_۾�k�����5	��]�!����M[��Ǣw�)��O�ҋX����>��l%i�-�M�g������{l�f|�ό���.���|��p��h�d �'���Xw�E�i�m}6*�3���f�]�!���D��L#�W�T ��x���� �+��T��/o��إP�e`b�T=am���� F����ȻD�ou�*Y x�S��q�©�����<�������~s���^��l8������t�iZ]XF��������;-;*�7��RTW�������&��J�1�KB|1<\w¹��<d�k�c��`��Z�>)��p40�zɈT^�`T�W�88�;矷A( ����_�h3��{I�B�+�7m_T���Q��K�����JU<o^.K�}��HwL�X'<�-Oɳ����=�Ҹ��H���~q4];ˍH��Σ"�]s=g����*F}Eo^��Ŏ>s��Y�&7�ܥ��2��
[���p�� +@���a
��|���\G�Y�)��Y�%�<'L�<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9���[�t��#����Ea��Z鎬�������(���P����ˮ��lC��U�T�\ ��+�_0c �X�FJ�+���-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0(����!
%Z鎬�������(���`$�P.eE���lC��U�T�\ ��+�_0c �w�)��O�ҋX����>��l%i�-�M�g������{l�f|�ό���.ӳ�
�	?�<7Ê7�E�4'���XwI<��f��F����U��:9�+�m��+���J q�v����6��w�1����R$b��m�+��
J��@��ea�8��������?9�f�*ʝ��%�}< V��,��B	hI�ˋ��b�ӝ5�T�@���k�փ��㛋��X���`��.�̀�I7��-5?�1J&�|D�e�!���QI�D/����ʊv.s/�B{�o
�Y-�E�f�}�=Ll�����,۽���}i�@�5�}�]���x�]�V��7��_��T��!e����\G�Y�)��Y櫧�7*9uu"�,�>E��<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9���[�t��#���j;9ekN�By3��<Z鎬�������(���P����ˮ��lC��U�T�\ ��+�_0c �Q�P��
S��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+�����
L'���Xw�j�7��ct�:��RE��W��_�ړ8���/�z&v��\��t������S�)37J*u>����C�/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�ЂDa��(O�J,���Z鎬����F�71�B��O1��m<S�)37J*u�񁫴}2;9�".<�x���� �+��T����oGo�Z�������--�p�,X�
���nx���� �+��T����oGo�Z�K����ހ d����f��WjCt�z&��ÃlO ܅dh�' L� U��֜��3jݭ�F���L�D��6S�]V�H7'�R�^Ƒ���a�\����9�	��%т��!o.sG[�� �`�>:8�A�/����<.+6J!�t���\�W��F�eD4];ˍH�7��_��T��!e����\G�YIpsl�ć���vh�ҋX������S8�J�]=��R�^Ƒ����"X��[��Q[R�7�%=��L�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y����q��G8�����b,�e.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7&�e��A�����
L'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<�e�y���J�@IE�U����S8�/ #O�)R�^Ƒ����"X��[�d�a�4$��9+�����o��C!T*�q���U����?�N�By3��<Z鎬�����X���*_��(֥�S�)37J*u>����CΫa������<��z��}���w�V�"-4��h�]8e�0
A���J��@��ea�8��������?9|[�,HJ
a�\7�"
qJH3#��Aq��:9�+�m��+�ڔ�wV��y�p�cP �����l8������t�iZ]XF�������� ��k\�\�KE���H���o��qo�:�ȓ��o)�]r k�|6�8��u*K6H.��h��u>j޽���Ǜ������[7�d|���XP��Ȩ�wl��h�Vx�%L��Ok��@zL͊�q���Vǃ���G&%	��ڔ��n����\�v�)��+�}��]�.�b�;װ?�p��U��֜��3JHn��z���G7�����o)�]rN�ǁ�f�T�J��H9��\�v�T?�7G|`^�R@Κ�2�Ix���KaJuA�����IÙ=�HF���m¡�3
�v�v-}�	mp�EN��S�IÙ=�H%v@����fnQ�rV4����X���\�v���GAџV^�R@Κ�2'�̗������\�ݠ�3zL͊�q��UG�s�����M���o�G�m�?M�*B�[zL͊�q��UG�s�����M���HaU$kX��� nU�IÙ=�HF���m¡A�h��+Fen����9��#�B�sYC��\�v��_�R�G�$����{v��G�K$xE�p4rqG7��u*K6H �i7�sp>��%��H��5[�����q�_�N�6�Ặ��Ϊ�Q� ~�����(��q�
�Bk�i�E?�xu����ma��u��ۯi\�q���Ì �&�k��>���c��d�|ݔ�3�5�}�]���x�]�V�����Ү��`�+S�p��ͷQ�X����fx'v�ao.\C�k�ף�D�~4#C(�}�IÙ=�H�%��@�Kǹ|���|u��RJHn��z��r9�3��X�u�ӑ�띂ii�4];ˍH���Vchw�D��y.���=��܄��띂ii�4];ˍH���Vchw�D��y.���eŞG�T(x�]�V���o��8���Cf֩Q�e]��W�'NTؕ@�.MŃ�,��)x�]�V���F�uB�W˪��/h�Б����x�]�V��,t����t�i�lK�I<��fҾ��9��ЂDa��(o��0��7��|g�Y�'���Xw�f�VHF��Q�#<4^�v�ј�"��Z鎬����F�71�B�������%�N�By3��<�]�!����M[��Ǣ�L ʞ��0��m��x���j���0z�cUL3�X�j��7$2Ӕ�1���_�wa(􆿳�tP"7��%e��0�U+�qbp@��wbk�$���7Z���(�
t�ژq���U� бb*	��|	�WI�����
L'���Xw�4��}�<�=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A����ɻ:�E�1N�By3��<�]�!���\B��V���#���L�
�����Yl���#�]�!��	Ǹ�y85��(�C)&���lC��U�T�\ �͹g}|�H���p��b��e������]�!��	Ǹ�y85���ǳ@�M�H�ɇM��lC��U�T�\ ��Tǯ�!���#;r�����S��I�?g�f��m���6d��h�Ɵ�Y�Ӿ���R$b�ȻD�ou�*Y x�S��q�©��L�=ɐ<c����4��G�p���ea�;y� ����t��o����q,� L��֍����A( ����_�h3��{I���s�ǘ5/��=��K��䘾is��E����F�'n�^0o��4�G�0�����Kp&�@���k��!�`�(i3�b9���j}8o{:�����Y�V�����ϲ������i��Q�^�y�zL͊�q���Vǃ���G&%	��ڏ�<
DN�!�`�(i3�b9���с�'sIP���1>y���Mw���1�Z���=��n̈́�zL͊�q��UG�s�����H(�T�O��{Tɀ���S�<Ԣ�JHn��z���o�K�Dd�KPZ���<om��������i�%Ah�%4
>��XP���nN#⦵���Օ��qvdЧ^{�j�E����F�'n�^0o��~+�ݗ�p�ϵ�DE1	�<�������Qt�2�b9����4�6�t�{]��ˀ.�� ��'���S ���3�ҺIÙ=�H��'�PD���ߜ�2a\c0@Ɓ��"�,�>E��ʆ�In��t�_�R�GI�~�џ0I� X�1�!�`�(i3���D	��U�l>o��|�w��Y�ڪ,[�=·j�C��[���Ԟ�����i����D	��U�l>o��|�w��Y�ڪ���E_����+�+#B�0|]<w:����D	��U�l>o��|���;�ĸ���_�?�)>*�7`����\Z��K���b9����4�6�t�g.��,��ҨԺ"�ߣ�g����=x�]�V�� �Gk	�}���f������r'��`m�oAr'�������i����D	��U�l>o��|��v���?�5�h�I�nI2z����!Cu�>(���] 9�Ln��S�W �i7�sp><F� ����/K��(�������i{!�`�(i3>���'hZ���j�Q%��{S'��{,�
w��|ݔ�3�(n�'��b9���:&�>��sw�n���7[q�m�J�5�d�,W�� nU�IÙ=�H��'�PD�A�h��+FeA'�u��o���T$�44];ˍH����Ү���/^�yQA�?��{m����
q<O�A'�u��o���T$�44];ˍH����Ү��`�+S�p��ͷQ�X��ފ�����x+�[Z��!�`�(i3x�]�V���	�?�ki%�7%1�e)s 3�:��)�[���6!�`�(i3���D	��U�l>o��|�,+$\�M��wF4��0[����	��N�Ae�#����ꀍ�����5	���]���>����C�h�'f RY%T��BPe.��xu	�>��l%i�-��9��稕�E����F��j��\w��0]ɍJ����j����tL��|g�Y�'���Xw�j�7��HaU$kX��a\Y���°��������ł�!r�dN�<@Iv��nt=:��(�
@��^y�~?�2vYl���#�]�!����M[��Ǣ+���G���"B��$I��w��,>����CΉ��S�|JY%T��BPe.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�� ߌ���E����F7G#+�Ǘ0z�cUL�BJ��VR�^Ƒ����"X��[��Q[R�7��=m緒��J���W�7G#+�Ǘ0z�cUL�J=��'EّD ����R�^Ƒ����"X��[�'i�! ]���f�e�0
A���J��@��ea�8���
ae���K�������
���nx���� �+��T���O'�lR�����|7!��CR��[ b�����,\ަ�ItK�1�֎TW������������i�l0��F��jT�����N��3w:��ݪ�򈟞�����i�%Ah�%4
>��XP������,��=�$�ЭU����z~��;ε��IÙ=�H:t@���8����̇i�d�?��E����F��j��\w��0]Y��
�iC"�,�>E����-��%Mό���.��6[��u�V�<�nbBIc��Et��q���U��X�=)�H�7M��񇬦���
L'���Xw��+x�r�2�6�d�f�]2�y�Z鎬����(��eظ�=�tneX N�By3��<�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+�� }'�8�������5	���]����,�JL���ƍ2���l�\.�l����"B��$I��w��,c�A�L'z��0N�7;�¬pX��g��U-�e�,���6+��kv޶Glbq�Z��T�I��w��,c�A�L'�b��9X�T��&��;�¬pX��g��U-�eaԗ5��C�Q�$�k\_x���� �+��T���O'�lR�����|7!��CR��U�
F�V�� VU+I��vMb��s��Yk"1/��n5R�%�.��.f\y㔪�_9&xc闑^����S����j�}�I/��=��K�R�/ؒ^�XzL͊�q����ϡ�����Kp&����-N���\�vņ�Q�]�ޔiyV�[R�^Ƒ���b9���j}8o{:��͹ ��1�Z���=�A ��E+���XP������,��=�$�ЭU����z~��;ε��IÙ=�HF���m¡�3
�v�v-}�	mp�EN��S�IÙ=�H�M�U�nQ�rV4����X���\�v�X�zgq��^�R@Κ�2'�̗������\�ݠ�3zL͊�q��UG�s�����M���o�G�m�?M�*B�[zL͊�q����![�_���S&ϊ�`�y���ʢȂ�zJ�^�R@Κ�2���C4�;��+���c�'n�^0o��~+�ݗ{,�
w��|ݔ�3�(n�'��b9���:&�>��sw�n���7[q�m�J�5�d�,W�� nU�IÙ=�H��'�PD�j�j2�%�5]��I踵}�=Ll�����&}0�@�͹ ��I�Q4p�/�;ϔW���1��ݥ�U� ���_�g)�X��Q�u������(�ʉ�I�,B�E?�xu����ma��u��ۯi\�q���Ìݣؤ	����2��̪C��[���ԍ�7�"�����=���aw��Y�ڪ,[�=·j�C��[���ԍ�7�"�����=���a��v6"S�����E_����+�+#B��1��ݥ�U� ���_?�(����ۙ��p�"�e|`����u�֗��}Eo^������m؅��FJ��������l�Y�f5/���i� � �	{����0�&�ͭ"�,�>E����-��%Mό���.��_F�k-�!�`�(i3c��Et��q���U��;���)"����}�����|g�Y�'���Xw�,bxqX��9��no��b�:/z��]���c�A�L'G~��6�7*���T��
����ѳ�T�\ �͘�f��p�b�z'hۉ)��d�7�q����B['u�E����F7G#+��\w��0]�r���h�0"�,�>E���TD��ό���.�q�\E��0M7$���c��Et�Y�{'%s��.|Z���I7��-5��6��	���`y�����sǪ��ɻ:�E�1N�By3��<�]�!���\B��V���q�-��H0�6GV�ꢤ�Og�[N�&ѐ�����
L'���Xw�j�7��U����z~��6��	���`y����*#�m z����Z��o�����
L'���Xw�j�7���=�$�ЭU����z~��6��	�\�HP@�a%=dϖ�i��F����U��:9�+�m��+�ڔ�wV���C�Sy6ג��̹��/R F����p�������.�<86�8m��+�����3�Χ��nEA�O����~